module top(in1, in2, in3, out1, out2);
input wire [15:0] in1;
input wire [15:0] in2;
input wire [15:0] in3;
output wire [31:0] out1;
output wire [31:0] out2;
assign w0 = ~in1[0];
assign w1 = ~in1[0];
assign w2 = ~in1[0];
assign w3 = ~in1[0];
assign w4 = ~in1[0];
assign w5 = ~in1[0];
assign w6 = in1[1] ~^ in1[0];
assign w7 = ~in1[1];
assign w8 = ~in1[1];
assign w9 = ~in1[1];
assign w10 = ~in1[1];
assign w11 = ~in1[1];
assign w12 = ~in1[1];
assign w13 = ~in1[1];
assign w14 = ~in1[1];
assign w15 = ~in1[1];
assign w16 = in1[2] ~^ in1[1];
assign w17 = ~in1[2];
assign w18 = ~in1[2];
assign w19 = ~in1[2];
assign w20 = ~in1[2];
assign w21 = ~in1[2];
assign w22 = ~in1[2];
assign w23 = ~in1[2];
assign w24 = ~in1[2];
assign w25 = ~in1[2];
assign w26 = in1[3] ~^ in1[2];
assign w27 = in1[3] ~| in1[2];
assign w28 = ~in1[3];
assign w29 = ~in1[3];
assign w30 = ~in1[3];
assign w31 = ~in1[3];
assign w32 = ~in1[3];
assign w33 = ~in1[3];
assign w34 = ~in1[3];
assign w35 = ~in1[3];
assign w36 = ~in1[3];
assign w37 = in1[4] ~^ in1[3];
assign w38 = in1[4] ~| in1[3];
assign w39 = ~in1[4];
assign w40 = ~in1[4];
assign w41 = ~in1[4];
assign w42 = ~in1[4];
assign w43 = ~in1[4];
assign w44 = ~in1[4];
assign w45 = ~in1[4];
assign w46 = ~in1[4];
assign w47 = ~in1[4];
assign w48 = in1[5] ~^ in1[4];
assign w49 = in1[5] ~| in1[4];
assign w50 = ~in1[5];
assign w51 = ~in1[5];
assign w52 = ~in1[5];
assign w53 = ~in1[5];
assign w54 = ~in1[5];
assign w55 = ~in1[5];
assign w56 = ~in1[5];
assign w57 = ~in1[5];
assign w58 = ~in1[5];
assign w59 = in1[6] ~^ in1[5];
assign w60 = in1[6] ~| in1[5];
assign w61 = ~in1[6];
assign w62 = ~in1[6];
assign w63 = ~in1[6];
assign w64 = ~in1[6];
assign w65 = ~in1[6];
assign w66 = ~in1[6];
assign w67 = ~in1[6];
assign w68 = ~in1[6];
assign w69 = ~in1[6];
assign w70 = in1[7] ~^ in1[6];
assign w71 = in1[7] ~| in1[6];
assign w72 = ~in1[7];
assign w73 = ~in1[7];
assign w74 = ~in1[7];
assign w75 = ~in1[7];
assign w76 = ~in1[7];
assign w77 = ~in1[7];
assign w78 = ~in1[7];
assign w79 = ~in1[7];
assign w80 = ~in1[7];
assign w81 = in1[8] ~^ in1[7];
assign w82 = in1[8] ~| in1[7];
assign w83 = ~in1[8];
assign w84 = ~in1[8];
assign w85 = ~in1[8];
assign w86 = ~in1[8];
assign w87 = ~in1[8];
assign w88 = ~in1[8];
assign w89 = ~in1[8];
assign w90 = ~in1[8];
assign w91 = ~in1[8];
assign w92 = in1[9] ~^ in1[8];
assign w93 = in1[9] ~| in1[8];
assign w94 = ~in1[9];
assign w95 = ~in1[9];
assign w96 = ~in1[9];
assign w97 = ~in1[9];
assign w98 = ~in1[9];
assign w99 = ~in1[9];
assign w100 = ~in1[9];
assign w101 = ~in1[9];
assign w102 = ~in1[9];
assign w103 = in1[10] ~^ in1[9];
assign w104 = in1[10] ~| in1[9];
assign w105 = ~in1[10];
assign w106 = ~in1[10];
assign w107 = ~in1[10];
assign w108 = ~in1[10];
assign w109 = ~in1[10];
assign w110 = ~in1[10];
assign w111 = ~in1[10];
assign w112 = ~in1[10];
assign w113 = ~in1[10];
assign w114 = in1[11] ~^ in1[10];
assign w115 = in1[11] ~| in1[10];
assign w116 = ~in1[11];
assign w117 = ~in1[11];
assign w118 = ~in1[11];
assign w119 = ~in1[11];
assign w120 = ~in1[11];
assign w121 = ~in1[11];
assign w122 = ~in1[11];
assign w123 = ~in1[11];
assign w124 = ~in1[11];
assign w125 = in1[12] ~^ in1[11];
assign w126 = in1[12] ~| in1[11];
assign w127 = ~in1[12];
assign w128 = ~in1[12];
assign w129 = ~in1[12];
assign w130 = ~in1[12];
assign w131 = ~in1[12];
assign w132 = ~in1[12];
assign w133 = ~in1[12];
assign w134 = ~in1[12];
assign w135 = ~in1[12];
assign w136 = in1[13] ~^ in1[12];
assign w137 = in1[13] ~| in1[12];
assign w138 = ~in1[13];
assign w139 = ~in1[13];
assign w140 = ~in1[13];
assign w141 = ~in1[13];
assign w142 = ~in1[13];
assign w143 = ~in1[13];
assign w144 = ~in1[13];
assign w145 = ~in1[13];
assign w146 = ~in1[13];
assign w147 = in1[14] ~^ in1[13];
assign w148 = in1[14] ~| in1[13];
assign w149 = ~in1[14];
assign w150 = ~in1[14];
assign w151 = ~in1[14];
assign w152 = ~in1[14];
assign w153 = ~in1[14];
assign w154 = ~in1[14];
assign w155 = ~in1[14];
assign w156 = ~in1[14];
assign w157 = ~in1[14];
assign w158 = in1[15] ~^ in1[14];
assign w159 = in1[15] ~| in1[14];
assign w160 = ~in1[15];
assign w161 = ~in1[15];
assign w162 = ~in1[15];
assign w163 = ~in1[15];
assign w164 = ~in1[15];
assign w165 = ~in1[15];
assign w166 = ~in1[15];
assign w167 = ~in1[15];
assign w168 = ~in1[15];
assign w169 = ~in2[0];
assign w170 = ~in2[1];
assign w171 = ~in2[2];
assign w172 = in2[3] ~^ in2[2];
assign w173 = ~in2[3];
assign w174 = ~in2[4];
assign w175 = ~in2[5];
assign w176 = in2[6] ~^ in2[5];
assign w177 = ~in2[6];
assign w178 = ~in2[7];
assign w179 = ~in2[8];
assign w180 = in2[9] ~^ in2[8];
assign w181 = ~in2[9];
assign w182 = ~in2[10];
assign w183 = ~in2[11];
assign w184 = in2[12] ~^ in2[11];
assign w185 = ~in2[12];
assign w186 = ~in2[13];
assign w187 = ~in2[14];
assign w188 = in2[15] & in2[14];
assign w189 = in2[15] ~| in2[14];
assign w190 = in2[2] | in3[0];
assign w191 = in2[2] & in3[0];
assign w192 = in2[5] ~^ in3[3];
assign w193 = in2[5] & in3[3];
assign w194 = in2[5] | in3[3];
assign w195 = in2[8] ~^ in3[6];
assign w196 = in2[8] | in3[6];
assign w197 = in2[8] & in3[6];
assign w198 = in2[11] ~^ in3[9];
assign w199 = in2[11] | in3[9];
assign w200 = in2[11] & in3[9];
assign w201 = in2[14] ~^ in3[12];
assign w202 = in2[14] | in3[12];
assign w203 = in2[14] & in3[12];
assign w204 = w3 | w7;
assign w205 = w12 | w25;
assign w206 = w17 | w30;
assign w207 = w28 | w44;
assign w208 = w39 | w50;
assign w209 = w55 | w61;
assign w210 = w66 | w77;
assign w211 = w72 | w83;
assign w212 = w88 | w99;
assign w213 = w94 | w105;
assign w214 = w110 | w121;
assign w215 = w116 | w127;
assign w216 = w132 | w143;
assign w217 = w138 | w154;
assign w218 = w149 | w168;
assign w219 = w170 | in2[0];
assign w220 = w171 ~^ in2[1];
assign w221 = w171 | in2[1];
assign w222 = w173 | in2[4];
assign w223 = w174 | in2[3];
assign w224 = in2[5] & w174;
assign w225 = w174 | in2[5];
assign w226 = w177 | in2[7];
assign w227 = w178 | in2[6];
assign w228 = in2[8] & w178;
assign w229 = w178 | in2[8];
assign w230 = w181 | in2[10];
assign w231 = w182 | in2[9];
assign w232 = in2[11] & w182;
assign w233 = w182 | in2[11];
assign w234 = w185 | in2[13];
assign w235 = w186 | in2[12];
assign w236 = in2[14] & w186;
assign w237 = w186 | in2[14];
assign w238 = ~w188;
assign w239 = ~w188;
assign w240 = ~w188;
assign w241 = ~w188;
assign w242 = ~w188;
assign w243 = ~w188;
assign w244 = ~w188;
assign w245 = ~w188;
assign w246 = w188 | w189;
assign w247 = w204 & w205;
assign w248 = w0 ~| w219;
assign w249 = w116 ~| w219;
assign w250 = w160 ~| w219;
assign w251 = w72 ~| w219;
assign w252 = w22 ~| w219;
assign w253 = w61 ~| w219;
assign w254 = w88 ~| w219;
assign w255 = w39 ~| w219;
assign w256 = w99 ~| w219;
assign w257 = w132 ~| w219;
assign w258 = w110 ~| w219;
assign w259 = w138 ~| w219;
assign w260 = w7 ~| w219;
assign w261 = w154 ~| w219;
assign w262 = w33 ~| w219;
assign w263 = w50 ~| w219;
assign w264 = w169 | w220;
assign w265 = ~w220;
assign w266 = in2[0] | w221;
assign w267 = w171 | w222;
assign w268 = in2[2] | w223;
assign w269 = ~w224;
assign w270 = w173 | w225;
assign w271 = ~w225;
assign w272 = w175 | w226;
assign w273 = in2[5] | w227;
assign w274 = ~w228;
assign w275 = w177 | w229;
assign w276 = ~w229;
assign w277 = w179 | w230;
assign w278 = in2[8] | w231;
assign w279 = ~w232;
assign w280 = w181 | w233;
assign w281 = ~w233;
assign w282 = w183 | w234;
assign w283 = in2[11] | w235;
assign w284 = ~w236;
assign w285 = w185 | w237;
assign w286 = ~w237;
assign w287 = w55 ~| w238;
assign w288 = w44 ~| w238;
assign w289 = w94 ~| w239;
assign w290 = w149 ~| w239;
assign w291 = w121 ~| w240;
assign w292 = w105 ~| w240;
assign w293 = w66 ~| w241;
assign w294 = w25 | w241;
assign w295 = w83 ~| w242;
assign w296 = w28 ~| w242;
assign w297 = w160 | w243;
assign w298 = w127 ~| w243;
assign w299 = w2 ~| w244;
assign w300 = w143 ~| w244;
assign w301 = w12 ~| w245;
assign w302 = w77 ~| w245;
assign w303 = w33 | w246;
assign w304 = ~w246;
assign w305 = ~w246;
assign w306 = ~w246;
assign w307 = ~w246;
assign w308 = ~w246;
assign w309 = ~w246;
assign w310 = ~w246;
assign w311 = ~w246;
assign w312 = w26 ~^ w247;
assign w313 = w27 | w247;
assign w314 = w11 ~| w264;
assign w315 = w43 ~| w264;
assign w316 = w119 ~| w264;
assign w317 = w98 ~| w264;
assign w318 = w109 ~| w264;
assign w319 = w153 ~| w264;
assign w320 = w84 ~| w264;
assign w321 = w54 ~| w264;
assign w322 = w165 ~| w264;
assign w323 = w142 ~| w264;
assign w324 = w32 ~| w264;
assign w325 = w18 ~| w264;
assign w326 = w76 ~| w264;
assign w327 = w131 ~| w264;
assign w328 = w64 ~| w264;
assign w329 = w169 | w265;
assign w330 = w96 ~| w266;
assign w331 = w1 ~| w266;
assign w332 = w107 ~| w266;
assign w333 = w74 ~| w266;
assign w334 = w129 ~| w266;
assign w335 = w9 ~| w266;
assign w336 = w19 ~| w266;
assign w337 = w140 ~| w266;
assign w338 = w85 ~| w266;
assign w339 = w151 ~| w266;
assign w340 = w165 ~| w266;
assign w341 = w52 ~| w266;
assign w342 = w63 ~| w266;
assign w343 = w41 ~| w266;
assign w344 = w118 ~| w266;
assign w345 = w35 ~| w266;
assign w346 = w267 & w268;
assign w347 = in2[3] ~| w269;
assign w348 = w171 ~| w270;
assign w349 = w224 | w271;
assign w350 = w272 & w273;
assign w351 = in2[6] ~| w274;
assign w352 = w175 ~| w275;
assign w353 = w228 | w276;
assign w354 = w277 & w278;
assign w355 = in2[9] ~| w279;
assign w356 = w179 ~| w280;
assign w357 = w232 | w281;
assign w358 = w282 & w283;
assign w359 = in2[12] ~| w284;
assign w360 = w183 ~| w285;
assign w361 = w236 | w286;
assign w362 = w294 & w303;
assign w363 = in1[11] & w304;
assign w364 = in1[12] & w304;
assign w365 = in1[15] & w305;
assign w366 = in1[7] & w305;
assign w367 = in1[8] & w306;
assign w368 = in1[5] & w306;
assign w369 = in1[0] & w307;
assign w370 = in1[1] & w307;
assign w371 = in1[2] & w308;
assign w372 = in1[14] & w308;
assign w373 = in1[13] & w309;
assign w374 = in1[9] & w309;
assign w375 = in1[6] & w310;
assign w376 = in1[4] & w310;
assign w377 = in1[10] & w311;
assign w378 = w206 & w313;
assign w379 = w312 ~| w329;
assign w380 = w264 & w329;
assign w381 = w6 ~| w329;
assign w382 = w258 | w330;
assign w383 = w260 | w331;
assign w384 = w249 | w332;
assign w385 = w254 | w333;
assign w386 = w259 | w334;
assign w387 = w252 | w335;
assign w388 = w262 | w336;
assign w389 = w261 | w337;
assign w390 = w256 | w338;
assign w391 = w250 | w339;
assign w392 = w253 | w341;
assign w393 = w251 | w342;
assign w394 = w263 | w343;
assign w395 = w257 | w344;
assign w396 = w255 | w345;
assign w397 = w0 ~| w346;
assign w398 = w30 ~| w346;
assign w399 = w162 ~| w346;
assign w400 = w119 ~| w346;
assign w401 = w39 ~| w346;
assign w402 = w20 ~| w346;
assign w403 = w64 ~| w346;
assign w404 = w130 ~| w346;
assign w405 = w14 ~| w346;
assign w406 = w51 ~| w346;
assign w407 = w79 ~| w346;
assign w408 = w101 ~| w346;
assign w409 = w86 ~| w346;
assign w410 = w152 ~| w346;
assign w411 = w108 ~| w346;
assign w412 = w141 ~| w346;
assign w413 = w171 & w347;
assign w414 = w172 | w349;
assign w415 = ~w349;
assign w416 = w5 ~| w350;
assign w417 = w86 ~| w350;
assign w418 = w10 ~| w350;
assign w419 = w65 ~| w350;
assign w420 = w53 ~| w350;
assign w421 = w97 ~| w350;
assign w422 = w152 ~| w350;
assign w423 = w130 ~| w350;
assign w424 = w72 ~| w350;
assign w425 = w123 ~| w350;
assign w426 = w46 ~| w350;
assign w427 = w145 ~| w350;
assign w428 = w166 ~| w350;
assign w429 = w30 ~| w350;
assign w430 = w17 ~| w350;
assign w431 = w112 ~| w350;
assign w432 = w175 & w351;
assign w433 = w176 | w353;
assign w434 = ~w353;
assign w435 = w4 ~| w354;
assign w436 = w97 ~| w354;
assign w437 = w161 ~| w354;
assign w438 = w108 ~| w354;
assign w439 = w42 ~| w354;
assign w440 = w73 ~| w354;
assign w441 = w53 ~| w354;
assign w442 = w68 ~| w354;
assign w443 = w8 ~| w354;
assign w444 = w139 ~| w354;
assign w445 = w150 ~| w354;
assign w446 = w117 ~| w354;
assign w447 = w28 ~| w354;
assign w448 = w90 ~| w354;
assign w449 = w20 ~| w354;
assign w450 = w128 ~| w354;
assign w451 = w179 & w355;
assign w452 = w180 | w357;
assign w453 = ~w357;
assign w454 = w1 ~| w358;
assign w455 = w62 ~| w358;
assign w456 = w163 ~| w358;
assign w457 = w120 ~| w358;
assign w458 = w22 ~| w358;
assign w459 = w95 ~| w358;
assign w460 = w87 ~| w358;
assign w461 = w156 ~| w358;
assign w462 = w75 ~| w358;
assign w463 = w141 ~| w358;
assign w464 = w42 ~| w358;
assign w465 = w57 ~| w358;
assign w466 = w10 ~| w358;
assign w467 = w134 ~| w358;
assign w468 = w106 ~| w358;
assign w469 = w29 ~| w358;
assign w470 = w183 & w359;
assign w471 = w184 | w361;
assign w472 = ~w361;
assign w473 = in2[2] | w362;
assign w474 = in2[2] & w362;
assign w475 = w292 | w363;
assign w476 = w291 | w364;
assign w477 = w290 | w365;
assign w478 = w293 | w366;
assign w479 = w302 | w367;
assign w480 = w288 | w368;
assign w481 = in3[15] & w369;
assign w482 = w369 ^ in3[15];
assign w483 = w299 | w370;
assign w484 = w301 | w371;
assign w485 = w300 | w372;
assign w486 = w298 | w373;
assign w487 = w295 | w374;
assign w488 = w287 | w375;
assign w489 = w296 | w376;
assign w490 = w289 | w377;
assign w491 = w37 ~^ w378;
assign w492 = w38 | w378;
assign w493 = w324 | w379;
assign w494 = w3 | w380;
assign w495 = w248 | w381;
assign w496 = w348 | w413;
assign w497 = w107 ~| w414;
assign w498 = w144 ~| w414;
assign w499 = w118 ~| w414;
assign w500 = w23 ~| w414;
assign w501 = w162 ~| w414;
assign w502 = w35 ~| w414;
assign w503 = w100 ~| w414;
assign w504 = w63 ~| w414;
assign w505 = w9 ~| w414;
assign w506 = w41 ~| w414;
assign w507 = w56 ~| w414;
assign w508 = w155 ~| w414;
assign w509 = w79 ~| w414;
assign w510 = w85 ~| w414;
assign w511 = w133 ~| w414;
assign w512 = w172 | w415;
assign w513 = w352 | w432;
assign w514 = w164 ~| w433;
assign w515 = w90 ~| w433;
assign w516 = w145 ~| w433;
assign w517 = w7 ~| w433;
assign w518 = w34 ~| w433;
assign w519 = w116 ~| w433;
assign w520 = w149 ~| w433;
assign w521 = w94 ~| w433;
assign w522 = w134 ~| w433;
assign w523 = w23 ~| w433;
assign w524 = w78 ~| w433;
assign w525 = w40 ~| w433;
assign w526 = w52 ~| w433;
assign w527 = w105 ~| w433;
assign w528 = w68 ~| w433;
assign w529 = w176 | w434;
assign w530 = w356 | w451;
assign w531 = w122 ~| w452;
assign w532 = w138 ~| w452;
assign w533 = w83 ~| w452;
assign w534 = w45 ~| w452;
assign w535 = w156 ~| w452;
assign w536 = w101 ~| w452;
assign w537 = w57 ~| w452;
assign w538 = w163 ~| w452;
assign w539 = w29 ~| w452;
assign w540 = w75 ~| w452;
assign w541 = w127 ~| w452;
assign w542 = w21 ~| w452;
assign w543 = w112 ~| w452;
assign w544 = w61 ~| w452;
assign w545 = w14 ~| w452;
assign w546 = w180 | w453;
assign w547 = w360 | w470;
assign w548 = w19 ~| w471;
assign w549 = w67 ~| w471;
assign w550 = w129 ~| w471;
assign w551 = w111 ~| w471;
assign w552 = w46 ~| w471;
assign w553 = w140 ~| w471;
assign w554 = w160 ~| w471;
assign w555 = w151 ~| w471;
assign w556 = w13 ~| w471;
assign w557 = w50 ~| w471;
assign w558 = w89 ~| w471;
assign w559 = w74 ~| w471;
assign w560 = w96 ~| w471;
assign w561 = w31 ~| w471;
assign w562 = w123 ~| w471;
assign w563 = w184 | w472;
assign w564 = ~w474;
assign w565 = ~w475;
assign w566 = w183 | w475;
assign w567 = w476 ~^ in2[11];
assign w568 = w477 ~^ in2[14];
assign w569 = ~w478;
assign w570 = ~w479;
assign w571 = w179 & w479;
assign w572 = ~w480;
assign w573 = w175 | w480;
assign w574 = w481 & w483;
assign w575 = w481 ^ w483;
assign w576 = ~w485;
assign w577 = w485 ~^ w486;
assign w578 = w187 | w486;
assign w579 = w487 ~^ in2[8];
assign w580 = w488 ~^ in2[5];
assign w581 = w474 ~| w489;
assign w582 = w474 ~^ w489;
assign w583 = ~w489;
assign w584 = ~w490;
assign w585 = w329 ~| w491;
assign w586 = w207 & w492;
assign w587 = w387 ~| w493;
assign w588 = w494 ~^ in2[2];
assign w589 = w314 ~| w495;
assign w590 = ~w496;
assign w591 = ~w496;
assign w592 = ~w496;
assign w593 = ~w496;
assign w594 = ~w496;
assign w595 = in1[0] & w496;
assign w596 = ~w496;
assign w597 = ~w496;
assign w598 = w405 | w500;
assign w599 = w410 | w501;
assign w600 = w409 | w503;
assign w601 = w401 | w507;
assign w602 = w412 | w508;
assign w603 = w407 | w510;
assign w604 = w312 ~| w512;
assign w605 = w414 & w512;
assign w606 = w491 ~| w512;
assign w607 = w6 ~| w512;
assign w608 = ~w513;
assign w609 = ~w513;
assign w610 = ~w513;
assign w611 = ~w513;
assign w612 = ~w513;
assign w613 = in1[0] & w513;
assign w614 = ~w513;
assign w615 = ~w513;
assign w616 = w431 | w519;
assign w617 = w417 | w521;
assign w618 = w425 | w522;
assign w619 = w421 | w527;
assign w620 = w312 ~| w529;
assign w621 = w433 & w529;
assign w622 = w491 ~| w529;
assign w623 = w6 ~| w529;
assign w624 = ~w530;
assign w625 = ~w530;
assign w626 = ~w530;
assign w627 = ~w530;
assign w628 = ~w530;
assign w629 = in1[0] & w530;
assign w630 = ~w530;
assign w631 = ~w530;
assign w632 = w440 | w533;
assign w633 = w447 | w534;
assign w634 = w439 | w537;
assign w635 = w449 | w539;
assign w636 = w442 | w540;
assign w637 = w446 | w541;
assign w638 = w443 | w542;
assign w639 = w441 | w544;
assign w640 = w435 | w545;
assign w641 = ~w546;
assign w642 = w491 ~| w546;
assign w643 = w6 ~| w546;
assign w644 = ~w547;
assign w645 = ~w547;
assign w646 = ~w547;
assign w647 = ~w547;
assign w648 = ~w547;
assign w649 = in1[0] & w547;
assign w650 = ~w547;
assign w651 = ~w547;
assign w652 = w466 | w548;
assign w653 = w465 | w549;
assign w654 = w469 | w552;
assign w655 = w454 | w556;
assign w656 = w464 | w557;
assign w657 = w458 | w561;
assign w658 = w468 | w562;
assign w659 = w312 ~| w563;
assign w660 = w471 & w563;
assign w661 = w491 ~| w563;
assign w662 = w6 ~| w563;
assign w663 = w473 & w564;
assign w664 = w490 | w565;
assign w665 = ~w565;
assign w666 = w476 & w566;
assign w667 = w475 ~^ w567;
assign w668 = w479 ~| w569;
assign w669 = w478 | w570;
assign w670 = ~w570;
assign w671 = w489 | w572;
assign w672 = ~w572;
assign w673 = w488 & w573;
assign w674 = w484 & w574;
assign w675 = w484 ^ w574;
assign w676 = w486 | w576;
assign w677 = w477 & w578;
assign w678 = w479 ~^ w579;
assign w679 = w480 ~^ w580;
assign w680 = w564 | w583;
assign w681 = w480 ~| w583;
assign w682 = w475 ~| w584;
assign w683 = w315 | w585;
assign w684 = w48 ~^ w586;
assign w685 = w49 | w586;
assign w686 = w587 ~^ in2[2];
assign w687 = w588 ~^ in2[2];
assign w688 = w190 & w588;
assign w689 = w589 ~^ in2[2];
assign w690 = w54 ~| w590;
assign w691 = w69 ~| w590;
assign w692 = w73 ~| w590;
assign w693 = w166 ~| w591;
assign w694 = w36 ~| w591;
assign w695 = w11 ~| w592;
assign w696 = w98 ~| w592;
assign w697 = w109 ~| w593;
assign w698 = w91 ~| w593;
assign w699 = w157 ~| w594;
assign w700 = w47 ~| w594;
assign w701 = w142 ~| w596;
assign w702 = w131 ~| w596;
assign w703 = w17 ~| w597;
assign w704 = w124 ~| w597;
assign w705 = w502 | w604;
assign w706 = w1 | w605;
assign w707 = w398 | w606;
assign w708 = w397 | w607;
assign w709 = w153 ~| w608;
assign w710 = w58 ~| w608;
assign w711 = w84 ~| w608;
assign w712 = w15 ~| w609;
assign w713 = w120 ~| w609;
assign w714 = w167 ~| w610;
assign w715 = w95 ~| w610;
assign w716 = w69 ~| w611;
assign w717 = w43 ~| w611;
assign w718 = w135 ~| w612;
assign w719 = w106 ~| w612;
assign w720 = w418 | w613;
assign w721 = w80 ~| w614;
assign w722 = w36 ~| w614;
assign w723 = w146 ~| w615;
assign w724 = w18 ~| w615;
assign w725 = w518 | w620;
assign w726 = w4 | w621;
assign w727 = w525 | w622;
assign w728 = w416 | w623;
assign w729 = w51 ~| w624;
assign w730 = w80 ~| w624;
assign w731 = w32 ~| w624;
assign w732 = w8 ~| w625;
assign w733 = w62 ~| w625;
assign w734 = w164 ~| w626;
assign w735 = w117 ~| w626;
assign w736 = w113 ~| w627;
assign w737 = w102 ~| w627;
assign w738 = w21 ~| w628;
assign w739 = w47 ~| w628;
assign w740 = w91 ~| w630;
assign w741 = w135 ~| w630;
assign w742 = w146 ~| w631;
assign w743 = w150 ~| w631;
assign w744 = ~w641;
assign w745 = w640 ~| w643;
assign w746 = w128 ~| w644;
assign w747 = w24 ~| w644;
assign w748 = w139 ~| w644;
assign w749 = w31 ~| w645;
assign w750 = w40 ~| w645;
assign w751 = w161 ~| w646;
assign w752 = w65 ~| w646;
assign w753 = w113 ~| w647;
assign w754 = w87 ~| w647;
assign w755 = w124 ~| w648;
assign w756 = w157 ~| w648;
assign w757 = w58 ~| w650;
assign w758 = w102 ~| w650;
assign w759 = w15 ~| w651;
assign w760 = w76 ~| w651;
assign w761 = w2 | w660;
assign w762 = w655 ~| w662;
assign w763 = ~w663;
assign w764 = w490 ~^ w665;
assign w765 = w183 & w665;
assign w766 = ~w667;
assign w767 = w478 ~^ w670;
assign w768 = w179 | w670;
assign w769 = w489 ~^ w672;
assign w770 = w175 & w672;
assign w771 = ~w674;
assign w772 = ~w678;
assign w773 = ~w679;
assign w774 = w388 ~| w683;
assign w775 = w329 ~| w684;
assign w776 = w546 ~| w684;
assign w777 = w563 ~| w684;
assign w778 = w512 ~| w684;
assign w779 = w529 ~| w684;
assign w780 = w208 & w685;
assign w781 = w687 ~^ in3[0];
assign w782 = w191 | w688;
assign w783 = w689 ~^ in3[1];
assign w784 = in3[1] & w689;
assign w785 = in3[1] | w689;
assign w786 = w403 | w690;
assign w787 = w402 | w695;
assign w788 = w411 | w696;
assign w789 = w400 | w697;
assign w790 = w408 | w698;
assign w791 = w399 | w699;
assign w792 = w406 | w700;
assign w793 = w506 | w703;
assign w794 = w404 | w704;
assign w795 = w706 ~^ in2[5];
assign w796 = w505 ~| w708;
assign w797 = w428 | w709;
assign w798 = w419 | w710;
assign w799 = w430 | w712;
assign w800 = w423 | w713;
assign w801 = w424 | w716;
assign w802 = w420 | w717;
assign w803 = w427 | w718;
assign w804 = w426 | w722;
assign w805 = w422 | w723;
assign w806 = w429 | w724;
assign w807 = w726 ~^ in2[8];
assign w808 = w517 ~| w728;
assign w809 = w448 | w730;
assign w810 = w532 | w735;
assign w811 = w438 | w737;
assign w812 = w642 | w738;
assign w813 = w436 | w740;
assign w814 = w444 | w741;
assign w815 = w445 | w742;
assign w816 = w437 | w743;
assign w817 = w312 ~| w744;
assign w818 = w452 & w744;
assign w819 = w745 ~^ in2[11];
assign w820 = w463 | w746;
assign w821 = w661 | w747;
assign w822 = w554 | w748;
assign w823 = w462 | w752;
assign w824 = w457 | w753;
assign w825 = w459 | w754;
assign w826 = w467 | w755;
assign w827 = w456 | w756;
assign w828 = w455 | w757;
assign w829 = w659 | w759;
assign w830 = w460 | w760;
assign w831 = w761 ~^ in2[14];
assign w832 = w762 ~^ in2[14];
assign w833 = w674 | w763;
assign w834 = w666 | w765;
assign w835 = w487 & w768;
assign w836 = w673 | w770;
assign w837 = w663 ~^ w771;
assign w838 = w663 ~| w771;
assign w839 = w774 ~^ in2[2];
assign w840 = w321 | w775;
assign w841 = w731 | w776;
assign w842 = w749 | w777;
assign w843 = w694 | w778;
assign w844 = w526 | w779;
assign w845 = w59 ~^ w780;
assign w846 = w60 | w780;
assign out2[0] = ~w781;
assign w847 = ~w781;
assign w848 = ~w781;
assign w849 = w782 ~^ w783;
assign w850 = w782 & w785;
assign w851 = w705 ~| w787;
assign w852 = w707 ~| w793;
assign w853 = w192 ~^ w795;
assign w854 = w194 & w795;
assign w855 = w796 ~^ in2[5];
assign w856 = w725 ~| w799;
assign w857 = w727 ~| w806;
assign w858 = w195 ~^ w807;
assign w859 = w196 & w807;
assign w860 = w808 ~^ in2[8];
assign w861 = w633 ~| w812;
assign w862 = w732 | w817;
assign w863 = w0 | w818;
assign w864 = w819 ~^ in3[10];
assign w865 = in3[10] | w819;
assign w866 = in3[10] & w819;
assign w867 = w654 ~| w821;
assign w868 = w657 ~| w829;
assign w869 = w201 ~^ w831;
assign w870 = w202 & w831;
assign w871 = w832 ~^ in3[13];
assign w872 = in3[13] | w832;
assign w873 = in3[13] & w832;
assign w874 = w486 ~^ w834;
assign w875 = w571 | w835;
assign w876 = w478 ~^ w836;
assign w877 = w569 & w836;
assign w878 = w569 | w836;
assign w879 = w396 ~| w840;
assign w880 = w634 ~| w841;
assign w881 = w656 ~| w842;
assign w882 = w601 ~| w843;
assign w883 = w804 ~| w844;
assign w884 = w512 ~| w845;
assign w885 = w563 ~| w845;
assign w886 = w329 ~| w845;
assign w887 = w546 ~| w845;
assign w888 = w529 ~| w845;
assign w889 = w209 & w846;
assign w890 = ~w848;
assign w891 = ~w849;
assign w892 = ~w849;
assign w893 = w784 | w850;
assign w894 = w851 ~^ in2[5];
assign w895 = w852 ~^ in2[5];
assign w896 = w686 ~^ w853;
assign w897 = w686 & w853;
assign w898 = w686 | w853;
assign w899 = w193 | w854;
assign w900 = in3[4] & w855;
assign w901 = in3[4] | w855;
assign w902 = w856 ~^ in2[8];
assign w903 = w857 ~^ in2[8];
assign w904 = w197 | w859;
assign w905 = w860 ~^ in3[7];
assign w906 = in3[7] & w860;
assign w907 = in3[7] | w860;
assign w908 = w861 ~^ in2[11];
assign w909 = w635 ~| w862;
assign w910 = w863 ~^ in2[11];
assign w911 = w867 ~^ in2[14];
assign w912 = w868 ~^ in2[14];
assign w913 = w203 | w870;
assign w914 = w490 ~^ w875;
assign w915 = w584 | w875;
assign w916 = w584 & w875;
assign w917 = w879 ~^ in2[2];
assign w918 = w880 ~^ in2[11];
assign w919 = w881 ~^ in2[14];
assign w920 = w882 ~^ in2[5];
assign w921 = w883 ~^ in2[8];
assign w922 = w504 | w884;
assign w923 = w750 | w885;
assign w924 = w328 | w886;
assign w925 = w739 | w887;
assign w926 = w528 | w888;
assign w927 = w70 ~^ w889;
assign w928 = w71 | w889;
assign w929 = w849 | w890;
assign w930 = w847 & w891;
assign w931 = w847 ~| w891;
assign w932 = w848 | w892;
assign w933 = w858 ~^ w894;
assign w934 = w858 | w894;
assign w935 = w858 & w894;
assign w936 = w899 ~^ in3[4];
assign w937 = w899 & w901;
assign w938 = w904 ~^ w905;
assign w939 = w904 & w907;
assign w940 = w909 ~^ in2[11];
assign w941 = w198 ~^ w910;
assign w942 = w199 & w910;
assign w943 = w575 ~^ w911;
assign w944 = w575 & w911;
assign w945 = w575 | w911;
assign w946 = w482 ~^ w912;
assign w947 = w482 & w912;
assign w948 = w482 | w912;
assign w949 = w871 ~^ w913;
assign w950 = w872 & w913;
assign w951 = w675 ~^ w919;
assign w952 = w675 & w919;
assign w953 = w675 | w919;
assign w954 = w792 ~| w922;
assign w955 = w653 ~| w923;
assign w956 = w394 ~| w924;
assign w957 = w639 ~| w925;
assign w958 = w802 ~| w926;
assign w959 = w563 ~| w927;
assign w960 = w529 ~| w927;
assign w961 = w546 ~| w927;
assign w962 = w512 ~| w927;
assign w963 = w329 ~| w927;
assign w964 = w210 & w928;
assign w965 = ~w930;
assign out2[1] = w930 | w931;
assign out1[1] = w929 & w932;
assign w966 = w855 ~^ w936;
assign w967 = w900 | w937;
assign w968 = w895 ~^ w938;
assign w969 = w895 | w938;
assign w970 = w895 & w938;
assign w971 = w906 | w939;
assign w972 = w869 ~^ w940;
assign w973 = w869 & w940;
assign w974 = w869 | w940;
assign w975 = w902 ~^ w941;
assign w976 = w902 & w941;
assign w977 = w902 | w941;
assign w978 = w200 | w942;
assign w979 = w908 ~^ w949;
assign w980 = w908 & w949;
assign w981 = w908 | w949;
assign w982 = w873 | w950;
assign w983 = w954 ~^ in2[5];
assign w984 = w955 ~^ in2[14];
assign w985 = w956 ~^ in2[2];
assign w986 = w957 ~^ in2[11];
assign w987 = w958 ~^ in2[8];
assign w988 = w559 | w959;
assign w989 = w524 | w960;
assign w990 = w729 | w961;
assign w991 = w509 | w962;
assign w992 = w326 | w963;
assign w993 = w81 ~^ w964;
assign w994 = w82 | w964;
assign w995 = w839 ~^ w966;
assign w996 = w839 | w966;
assign w997 = w839 & w966;
assign w998 = w864 ~^ w978;
assign w999 = w865 & w978;
assign w1000 = w837 ~^ w984;
assign w1001 = w833 & w984;
assign w1002 = w828 ~| w988;
assign w1003 = w798 ~| w989;
assign w1004 = w636 ~| w990;
assign w1005 = w786 ~| w991;
assign w1006 = w392 ~| w992;
assign w1007 = w512 ~| w993;
assign w1008 = w529 ~| w993;
assign w1009 = ~w993;
assign w1010 = w211 & w994;
assign w1011 = w903 ~^ w998;
assign w1012 = w903 & w998;
assign w1013 = w903 | w998;
assign w1014 = w866 | w999;
assign w1015 = w838 | w1001;
assign w1016 = w1002 ~^ in2[14];
assign w1017 = w1003 ~^ in2[8];
assign w1018 = w1004 ~^ in2[11];
assign w1019 = w1005 ~^ in2[5];
assign w1020 = w1006 ~^ in2[2];
assign w1021 = w691 | w1007;
assign w1022 = w515 | w1008;
assign w1023 = ~w1009;
assign w1024 = w641 & w1009;
assign w1025 = w92 ~^ w1010;
assign w1026 = w93 | w1010;
assign w1027 = w582 ~^ w1016;
assign w1028 = w680 & w1016;
assign w1029 = w603 ~| w1021;
assign w1030 = w801 ~| w1022;
assign w1031 = w329 ~| w1023;
assign w1032 = w563 ~| w1023;
assign w1033 = w733 | w1024;
assign w1034 = w546 ~| w1025;
assign w1035 = w563 ~| w1025;
assign w1036 = w329 ~| w1025;
assign w1037 = w529 ~| w1025;
assign w1038 = w512 ~| w1025;
assign w1039 = w212 & w1026;
assign w1040 = w1015 ~^ w1027;
assign w1041 = w1015 & w1027;
assign w1042 = w1015 | w1027;
assign w1043 = w581 | w1028;
assign w1044 = w1029 ~^ in2[5];
assign w1045 = w1030 ~^ in2[8];
assign w1046 = w320 | w1031;
assign w1047 = w558 | w1032;
assign w1048 = w632 ~| w1033;
assign w1049 = w536 | w1034;
assign w1050 = w560 | w1035;
assign w1051 = w317 | w1036;
assign w1052 = w721 | w1037;
assign w1053 = w692 | w1038;
assign w1054 = w103 ~^ w1039;
assign w1055 = w104 | w1039;
assign w1056 = ~w1043;
assign w1057 = w393 ~| w1046;
assign w1058 = w823 ~| w1047;
assign w1059 = w1048 ~^ in2[11];
assign w1060 = w809 ~| w1049;
assign w1061 = w830 ~| w1050;
assign w1062 = w385 ~| w1051;
assign w1063 = w617 ~| w1052;
assign w1064 = w600 ~| w1053;
assign w1065 = w563 ~| w1054;
assign w1066 = w529 ~| w1054;
assign w1067 = w329 ~| w1054;
assign w1068 = w546 ~| w1054;
assign w1069 = w512 ~| w1054;
assign w1070 = w213 & w1055;
assign w1071 = w1057 ~^ in2[2];
assign w1072 = w1058 ~^ in2[14];
assign w1073 = w1060 ~^ in2[11];
assign w1074 = w1061 ~^ in2[14];
assign w1075 = w1062 ~^ in2[2];
assign w1076 = w1063 ~^ in2[8];
assign w1077 = w1064 ~^ in2[5];
assign w1078 = w551 | w1065;
assign w1079 = w711 | w1066;
assign w1080 = w318 | w1067;
assign w1081 = w543 | w1068;
assign w1082 = w497 | w1069;
assign w1083 = w114 ~^ w1070;
assign w1084 = w115 | w1070;
assign w1085 = w769 ~^ w1072;
assign w1086 = w671 & w1072;
assign w1087 = w679 ~^ w1074;
assign w1088 = w773 | w1074;
assign w1089 = ~w1074;
assign w1090 = w825 ~| w1078;
assign w1091 = w619 ~| w1079;
assign w1092 = w390 ~| w1080;
assign w1093 = w813 ~| w1081;
assign w1094 = w790 ~| w1082;
assign w1095 = w512 ~| w1083;
assign w1096 = w563 ~| w1083;
assign w1097 = w329 ~| w1083;
assign w1098 = w546 ~| w1083;
assign w1099 = w529 ~| w1083;
assign w1100 = w214 & w1084;
assign w1101 = w1043 ~^ w1085;
assign w1102 = w1056 ~| w1085;
assign w1103 = ~w1085;
assign w1104 = w681 | w1086;
assign w1105 = w679 ~| w1089;
assign w1106 = w1090 ~^ in2[14];
assign w1107 = w1091 ~^ in2[8];
assign w1108 = w1092 ~^ in2[2];
assign w1109 = w1093 ~^ in2[11];
assign w1110 = w1094 ~^ in2[5];
assign w1111 = w499 | w1095;
assign w1112 = w758 | w1096;
assign w1113 = w316 | w1097;
assign w1114 = w531 | w1098;
assign w1115 = w715 | w1099;
assign w1116 = w125 ~^ w1100;
assign w1117 = w126 | w1100;
assign w1118 = w1043 | w1103;
assign w1119 = w1087 ~^ w1104;
assign w1120 = w1088 & w1104;
assign w1121 = w876 ~^ w1106;
assign w1122 = w878 & w1106;
assign w1123 = w1040 ~^ w1109;
assign w1124 = w1042 & w1109;
assign w1125 = w788 ~| w1111;
assign w1126 = w658 ~| w1112;
assign w1127 = w382 ~| w1113;
assign w1128 = w811 ~| w1114;
assign w1129 = w616 ~| w1115;
assign w1130 = w512 ~| w1116;
assign w1131 = w563 ~| w1116;
assign w1132 = w546 ~| w1116;
assign w1133 = w329 ~| w1116;
assign w1134 = w529 ~| w1116;
assign w1135 = w215 & w1117;
assign w1136 = ~w1119;
assign w1137 = w1105 | w1120;
assign w1138 = ~w1121;
assign w1139 = w877 | w1122;
assign w1140 = w1041 | w1124;
assign w1141 = w1125 ~^ in2[5];
assign w1142 = w1126 ~^ in2[14];
assign w1143 = w1127 ~^ in2[2];
assign w1144 = w1128 ~^ in2[11];
assign w1145 = w1129 ~^ in2[8];
assign w1146 = w511 | w1130;
assign w1147 = w550 | w1131;
assign w1148 = w736 | w1132;
assign w1149 = w327 | w1133;
assign w1150 = w719 | w1134;
assign w1151 = w136 ~^ w1135;
assign w1152 = w137 | w1135;
assign w1153 = w1121 ~^ w1137;
assign w1154 = ~w1137;
assign w1155 = w1137 | w1138;
assign w1156 = ~w1139;
assign w1157 = ~w1140;
assign w1158 = w767 ~^ w1142;
assign w1159 = w669 & w1142;
assign w1160 = w1101 ~^ w1144;
assign w1161 = w1118 & w1144;
assign w1162 = w789 ~| w1146;
assign w1163 = w824 ~| w1147;
assign w1164 = w637 ~| w1148;
assign w1165 = w384 ~| w1149;
assign w1166 = w618 ~| w1150;
assign w1167 = w329 ~| w1151;
assign w1168 = w563 ~| w1151;
assign w1169 = w512 ~| w1151;
assign w1170 = w529 ~| w1151;
assign w1171 = w546 ~| w1151;
assign w1172 = w216 & w1152;
assign w1173 = w1121 ~| w1154;
assign w1174 = w1139 ~^ w1158;
assign w1175 = w1156 ~| w1158;
assign w1176 = ~w1158;
assign w1177 = w668 | w1159;
assign w1178 = w1140 ~^ w1160;
assign w1179 = w1157 ~| w1160;
assign w1180 = ~w1160;
assign w1181 = w1102 | w1161;
assign w1182 = w1162 ~^ in2[5];
assign w1183 = w1163 ~^ in2[14];
assign w1184 = w1164 ~^ in2[11];
assign w1185 = w1165 ~^ in2[2];
assign w1186 = w1166 ~^ in2[8];
assign w1187 = w323 | w1167;
assign w1188 = w553 | w1168;
assign w1189 = w498 | w1169;
assign w1190 = w516 | w1170;
assign w1191 = w450 | w1171;
assign w1192 = w147 ~^ w1172;
assign w1193 = w148 | w1172;
assign w1194 = w1139 | w1176;
assign w1195 = w1140 | w1180;
assign w1196 = w678 ~^ w1183;
assign w1197 = w772 | w1183;
assign w1198 = ~w1183;
assign w1199 = w1119 ~^ w1184;
assign w1200 = w1136 | w1184;
assign w1201 = ~w1184;
assign w1202 = w395 ~| w1187;
assign w1203 = w826 ~| w1188;
assign w1204 = w794 ~| w1189;
assign w1205 = w800 ~| w1190;
assign w1206 = w810 ~| w1191;
assign w1207 = w529 ~| w1192;
assign w1208 = w329 ~| w1192;
assign w1209 = w563 ~| w1192;
assign w1210 = w512 ~| w1192;
assign w1211 = w546 ~| w1192;
assign w1212 = w217 & w1193;
assign w1213 = w1177 ~^ w1196;
assign w1214 = w1177 & w1197;
assign w1215 = w678 ~| w1198;
assign w1216 = w1181 ~^ w1199;
assign w1217 = w1181 & w1200;
assign w1218 = w1119 ~| w1201;
assign w1219 = w1202 ~^ in2[2];
assign w1220 = w1203 ~^ in2[14];
assign w1221 = w1204 ~^ in2[5];
assign w1222 = w1205 ~^ in2[8];
assign w1223 = w1206 ~^ in2[11];
assign w1224 = w520 | w1207;
assign w1225 = w319 | w1208;
assign w1226 = w555 | w1209;
assign w1227 = w702 | w1210;
assign w1228 = w535 | w1211;
assign w1229 = w158 ~^ w1212;
assign w1230 = w159 | w1212;
assign w1231 = ~w1213;
assign w1232 = w1214 | w1215;
assign w1233 = ~w1216;
assign w1234 = w1217 | w1218;
assign w1235 = w914 ~^ w1220;
assign w1236 = w915 & w1220;
assign w1237 = w1153 ~^ w1223;
assign w1238 = w1155 & w1223;
assign w1239 = w803 ~| w1224;
assign w1240 = w386 ~| w1225;
assign w1241 = w820 ~| w1226;
assign w1242 = w602 ~| w1227;
assign w1243 = w814 ~| w1228;
assign w1244 = w529 ~| w1229;
assign w1245 = w563 ~| w1229;
assign w1246 = w329 ~| w1229;
assign w1247 = w512 ~| w1229;
assign w1248 = w546 ~| w1229;
assign w1249 = w218 & w1230;
assign w1250 = ~w1232;
assign w1251 = ~w1234;
assign w1252 = w1232 ~^ w1235;
assign w1253 = ~w1235;
assign w1254 = w916 | w1236;
assign w1255 = w1234 ~^ w1237;
assign w1256 = ~w1237;
assign w1257 = w1173 | w1238;
assign w1258 = w1239 ~^ in2[8];
assign w1259 = w1240 ~^ in2[2];
assign w1260 = w1241 ~^ in2[14];
assign w1261 = w1242 ~^ in2[5];
assign w1262 = w1243 ~^ in2[11];
assign w1263 = w514 | w1244;
assign w1264 = w461 | w1245;
assign w1265 = w322 | w1246;
assign w1266 = w701 | w1247;
assign w1267 = w538 | w1248;
assign w1268 = w168 | w1249;
assign w1269 = ~w1249;
assign w1270 = w1235 ~| w1250;
assign w1271 = w1237 ~| w1251;
assign w1272 = w1232 | w1253;
assign w1273 = ~w1254;
assign w1274 = w1234 | w1256;
assign w1275 = ~w1257;
assign w1276 = w1178 ~^ w1258;
assign w1277 = w1195 & w1258;
assign w1278 = w764 ~^ w1260;
assign w1279 = w664 & w1260;
assign w1280 = w1174 ~^ w1262;
assign w1281 = w1194 & w1262;
assign w1282 = w805 ~| w1263;
assign w1283 = w822 ~| w1264;
assign w1284 = w389 ~| w1265;
assign w1285 = w599 ~| w1266;
assign w1286 = w815 ~| w1267;
assign w1287 = w529 ~| w1268;
assign w1288 = w546 ~| w1268;
assign w1289 = w563 ~| w1268;
assign w1290 = w512 ~| w1268;
assign w1291 = ~w1268;
assign w1292 = w329 ~| w1268;
assign w1293 = in1[15] ~| w1269;
assign w1294 = w1179 | w1277;
assign w1295 = w1254 ~^ w1278;
assign w1296 = w682 | w1279;
assign w1297 = w1257 ~^ w1280;
assign w1298 = w1175 | w1281;
assign w1299 = w1282 ~^ in2[8];
assign w1300 = w1283 ~^ in2[14];
assign w1301 = w1284 ~^ in2[2];
assign w1302 = w1285 ~^ in2[5];
assign w1303 = w1286 ~^ in2[11];
assign w1304 = w714 | w1287;
assign w1305 = w734 | w1288;
assign w1306 = w751 | w1289;
assign w1307 = w693 | w1290;
assign w1308 = w340 | w1292;
assign w1309 = w1291 | w1293;
assign w1310 = w1216 ~^ w1299;
assign w1311 = w1233 | w1299;
assign w1312 = ~w1299;
assign w1313 = w667 ~^ w1300;
assign w1314 = w766 | w1300;
assign w1315 = ~w1300;
assign w1316 = w1213 ~^ w1303;
assign w1317 = w1231 | w1303;
assign w1318 = ~w1303;
assign w1319 = w1304 ~^ in2[8];
assign w1320 = w1305 ~^ in2[11];
assign w1321 = w1306 ~^ in2[14];
assign w1322 = w1307 ~^ in2[5];
assign w1323 = w1308 ~^ in2[2];
assign w1324 = w329 ~| w1309;
assign w1325 = w529 ~| w1309;
assign w1326 = w512 ~| w1309;
assign w1327 = w546 ~| w1309;
assign w1328 = w563 ~| w1309;
assign w1329 = w1294 ~^ w1310;
assign w1330 = w1294 & w1311;
assign w1331 = w1216 ~| w1312;
assign w1332 = w1296 ~^ w1313;
assign w1333 = w1296 & w1314;
assign w1334 = w667 ~| w1315;
assign w1335 = w1298 ~^ w1316;
assign w1336 = w1298 & w1317;
assign w1337 = w1213 ~| w1318;
assign w1338 = w1297 ~^ w1319;
assign w1339 = w1275 | w1319;
assign w1340 = ~w1319;
assign w1341 = w1295 ~^ w1320;
assign w1342 = w1273 | w1320;
assign w1343 = ~w1320;
assign w1344 = w577 ~^ w1321;
assign w1345 = ~w1322;
assign w1346 = w391 ~| w1324;
assign w1347 = w797 ~| w1325;
assign w1348 = w791 ~| w1326;
assign w1349 = w816 ~| w1327;
assign w1350 = w827 ~| w1328;
assign w1351 = w1330 | w1331;
assign w1352 = w1333 | w1334;
assign w1353 = w1336 | w1337;
assign w1354 = w1257 ~| w1340;
assign w1355 = ~w1341;
assign w1356 = w1254 ~| w1343;
assign w1357 = w1346 ~^ in2[2];
assign w1358 = w1347 ~^ in2[8];
assign w1359 = w1348 ~^ in2[5];
assign w1360 = w1349 ~^ in2[11];
assign w1361 = w1350 ~^ in2[14];
assign w1362 = ~w1351;
assign w1363 = ~w1352;
assign w1364 = ~w1353;
assign w1365 = w1280 | w1354;
assign w1366 = w1278 | w1356;
assign w1367 = w1255 ~^ w1358;
assign w1368 = w1274 & w1358;
assign w1369 = w1252 ~^ w1360;
assign w1370 = w1272 & w1360;
assign w1371 = w874 ~^ w1361;
assign w1372 = w1339 & w1365;
assign w1373 = w1342 & w1366;
assign w1374 = w1351 ~^ w1367;
assign w1375 = w1362 ~| w1367;
assign w1376 = w1362 & w1367;
assign w1377 = w1271 | w1368;
assign w1378 = w1353 ~^ w1369;
assign w1379 = w1364 | w1369;
assign w1380 = ~w1369;
assign w1381 = w1270 | w1370;
assign w1382 = w1352 ~^ w1371;
assign w1383 = w1363 & w1371;
assign w1384 = w1363 ~| w1371;
assign w1385 = w1335 ~^ w1372;
assign w1386 = w1335 | w1372;
assign w1387 = w1335 & w1372;
assign w1388 = w1332 ~^ w1373;
assign w1389 = w1332 | w1373;
assign w1390 = w1332 & w1373;
assign w1391 = w1338 ~^ w1377;
assign w1392 = w1338 | w1377;
assign w1393 = w1338 & w1377;
assign w1394 = w1353 ~| w1380;
assign w1395 = w1341 ~^ w1381;
assign w1396 = w1341 ~| w1381;
assign w1397 = ~w1381;
assign w1398 = w1355 | w1397;
wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398;
endmodule
module top(in1, in2, in3, in4, in5, in6, out1, out2, out3, out4, out5);
input wire [1:0] in1;
input wire [1:0] in2;
input wire [4:0] in3;
input wire [2:0] in4;
input wire [4:0] in5;
input wire [2:0] in6;
output wire [4:0] out1;
output wire out2;
output wire [4:0] out3;
output wire out4;
output wire [4:0] out5;

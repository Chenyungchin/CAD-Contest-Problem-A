module top(in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, out1);
input wire [8:0] in1;
input wire in10;
input wire in11;
input wire [8:0] in12;
input wire [7:0] in13;
input wire in14;
input wire in15;
input wire [8:0] in16;
input wire [7:0] in17;
input wire in18;
input wire in19;
input wire [7:0] in2;
input wire [8:0] in20;
input wire [7:0] in21;
input wire in22;
input wire in23;
input wire [8:0] in24;
input wire [7:0] in25;
input wire in3;
input wire in4;
input wire [6:0] in5;
input wire in6;
input wire in7;
input wire [8:0] in8;
input wire [7:0] in9;
output wire [16:0] out1;
assign w0 = ~in10;
assign w1 = ~in10;
assign w2 = ~in12[0];
assign w3 = ~in12[1];
assign w4 = ~in12[2];
assign w5 = ~in12[3];
assign w6 = ~in12[4];
assign w7 = ~in12[5];
assign w8 = ~in12[6];
assign w9 = ~in12[7];
assign w10 = ~in12[8];
assign w11 = in12[5] & in13[0];
assign w12 = in12[3] & in13[0];
assign w13 = in12[4] & in13[0];
assign w14 = in12[6] & in13[0];
assign w15 = ~in13[0];
assign w16 = in12[8] & in13[1];
assign w17 = in12[4] & in13[1];
assign w18 = ~in13[1];
assign w19 = in12[7] & in13[2];
assign w20 = ~in13[2];
assign w21 = ~in13[3];
assign w22 = ~in13[4];
assign w23 = in12[3] & in13[5];
assign w24 = in12[0] & in13[5];
assign w25 = ~in13[5];
assign w26 = in12[2] & in13[6];
assign w27 = ~in13[6];
assign w28 = in12[8] & in13[7];
assign w29 = ~in13[7];
assign w30 = ~in14;
assign w31 = ~in14;
assign w32 = ~in16[0];
assign w33 = ~in16[1];
assign w34 = ~in16[2];
assign w35 = ~in16[3];
assign w36 = ~in16[4];
assign w37 = ~in16[5];
assign w38 = ~in16[6];
assign w39 = ~in16[7];
assign w40 = ~in16[8];
assign w41 = in16[5] & in17[0];
assign w42 = in16[3] & in17[0];
assign w43 = in16[4] & in17[0];
assign w44 = in16[6] & in17[0];
assign w45 = ~in17[0];
assign w46 = in16[8] & in17[1];
assign w47 = in16[4] & in17[1];
assign w48 = ~in17[1];
assign w49 = in16[7] & in17[2];
assign w50 = ~in17[2];
assign w51 = ~in17[3];
assign w52 = ~in17[4];
assign w53 = in16[3] & in17[5];
assign w54 = in16[0] & in17[5];
assign w55 = ~in17[5];
assign w56 = in16[2] & in17[6];
assign w57 = ~in17[6];
assign w58 = in16[8] & in17[7];
assign w59 = ~in17[7];
assign w60 = ~in18;
assign w61 = ~in18;
assign w62 = ~in1[0];
assign w63 = ~in1[1];
assign w64 = ~in1[2];
assign w65 = ~in1[3];
assign w66 = ~in1[4];
assign w67 = ~in1[5];
assign w68 = ~in1[6];
assign w69 = ~in1[7];
assign w70 = ~in1[8];
assign w71 = ~in20[0];
assign w72 = ~in20[1];
assign w73 = ~in20[2];
assign w74 = ~in20[3];
assign w75 = ~in20[4];
assign w76 = ~in20[5];
assign w77 = ~in20[6];
assign w78 = ~in20[7];
assign w79 = ~in20[8];
assign w80 = in20[5] & in21[0];
assign w81 = in20[3] & in21[0];
assign w82 = in20[4] & in21[0];
assign w83 = in20[6] & in21[0];
assign w84 = ~in21[0];
assign w85 = in20[8] & in21[1];
assign w86 = in20[4] & in21[1];
assign w87 = ~in21[1];
assign w88 = in20[7] & in21[2];
assign w89 = ~in21[2];
assign w90 = ~in21[3];
assign w91 = ~in21[4];
assign w92 = in20[3] & in21[5];
assign w93 = in20[0] & in21[5];
assign w94 = ~in21[5];
assign w95 = in20[2] & in21[6];
assign w96 = ~in21[6];
assign w97 = in20[8] & in21[7];
assign w98 = ~in21[7];
assign w99 = ~in22;
assign w100 = ~in22;
assign w101 = ~in24[0];
assign w102 = ~in24[1];
assign w103 = ~in24[2];
assign w104 = ~in24[3];
assign w105 = ~in24[4];
assign w106 = ~in24[5];
assign w107 = ~in24[6];
assign w108 = ~in24[7];
assign w109 = ~in24[8];
assign w110 = in24[5] & in25[0];
assign w111 = in24[3] & in25[0];
assign w112 = in24[4] & in25[0];
assign w113 = in24[6] & in25[0];
assign w114 = ~in25[0];
assign w115 = in24[8] & in25[1];
assign w116 = in24[4] & in25[1];
assign w117 = ~in25[1];
assign w118 = in24[7] & in25[2];
assign w119 = ~in25[2];
assign w120 = ~in25[3];
assign w121 = ~in25[4];
assign w122 = in24[3] & in25[5];
assign w123 = in24[0] & in25[5];
assign w124 = ~in25[5];
assign w125 = in24[2] & in25[6];
assign w126 = ~in25[6];
assign w127 = in24[8] & in25[7];
assign w128 = ~in25[7];
assign w129 = in1[5] & in2[0];
assign w130 = in1[3] & in2[0];
assign w131 = in1[4] & in2[0];
assign w132 = in1[6] & in2[0];
assign w133 = ~in2[0];
assign w134 = in1[8] & in2[1];
assign w135 = in1[4] & in2[1];
assign w136 = ~in2[1];
assign w137 = in1[7] & in2[2];
assign w138 = ~in2[2];
assign w139 = ~in2[3];
assign w140 = ~in2[4];
assign w141 = in1[3] & in2[5];
assign w142 = in1[0] & in2[5];
assign w143 = ~in2[5];
assign w144 = in1[2] & in2[6];
assign w145 = ~in2[6];
assign w146 = in1[8] & in2[7];
assign w147 = ~in2[7];
assign w148 = ~in3;
assign w149 = ~in3;
assign w150 = ~in5[1];
assign w151 = ~in5[2];
assign w152 = ~in5[3];
assign w153 = ~in6;
assign w154 = ~in6;
assign w155 = ~in8[0];
assign w156 = ~in8[1];
assign w157 = ~in8[2];
assign w158 = ~in8[3];
assign w159 = ~in8[4];
assign w160 = ~in8[5];
assign w161 = ~in8[6];
assign w162 = ~in8[7];
assign w163 = ~in8[8];
assign w164 = in8[5] & in9[0];
assign w165 = in8[3] & in9[0];
assign w166 = in8[4] & in9[0];
assign w167 = in8[6] & in9[0];
assign w168 = ~in9[0];
assign w169 = in8[8] & in9[1];
assign w170 = in8[4] & in9[1];
assign w171 = ~in9[1];
assign w172 = in8[7] & in9[2];
assign w173 = ~in9[2];
assign w174 = ~in9[3];
assign w175 = ~in9[4];
assign w176 = in8[3] & in9[5];
assign w177 = in8[0] & in9[5];
assign w178 = ~in9[5];
assign w179 = in8[2] & in9[6];
assign w180 = ~in9[6];
assign w181 = in8[8] & in9[7];
assign w182 = ~in9[7];
assign w183 = ~w0;
assign w184 = ~w1;
assign w185 = ~w2;
assign w186 = ~w2;
assign w187 = ~w3;
assign w188 = ~w3;
assign w189 = ~w4;
assign w190 = ~w4;
assign w191 = ~w5;
assign w192 = ~w5;
assign w193 = ~w6;
assign w194 = ~w6;
assign w195 = ~w7;
assign w196 = ~w7;
assign w197 = ~w8;
assign w198 = ~w8;
assign w199 = ~w9;
assign w200 = ~w9;
assign w201 = ~w10;
assign w202 = ~w10;
assign w203 = ~w15;
assign w204 = w11 & w17;
assign w205 = w11 ~^ w17;
assign w206 = ~w18;
assign w207 = w16 & w19;
assign w208 = w16 ~^ w19;
assign w209 = ~w20;
assign w210 = ~w20;
assign w211 = ~w21;
assign w212 = ~w21;
assign w213 = ~w21;
assign w214 = ~w22;
assign w215 = ~w22;
assign w216 = ~w22;
assign w217 = ~w23;
assign w218 = ~w24;
assign w219 = ~w25;
assign w220 = ~w25;
assign w221 = w23 | w26;
assign w222 = ~w26;
assign w223 = ~w27;
assign w224 = ~w27;
assign w225 = ~w29;
assign w226 = ~w29;
assign w227 = ~w30;
assign w228 = ~w31;
assign w229 = ~w32;
assign w230 = ~w32;
assign w231 = ~w33;
assign w232 = ~w33;
assign w233 = ~w34;
assign w234 = ~w34;
assign w235 = ~w35;
assign w236 = ~w35;
assign w237 = ~w36;
assign w238 = ~w36;
assign w239 = ~w37;
assign w240 = ~w37;
assign w241 = ~w38;
assign w242 = ~w38;
assign w243 = ~w39;
assign w244 = ~w39;
assign w245 = ~w40;
assign w246 = ~w40;
assign w247 = ~w45;
assign w248 = w41 & w47;
assign w249 = w41 ~^ w47;
assign w250 = ~w48;
assign w251 = w46 & w49;
assign w252 = w46 ~^ w49;
assign w253 = ~w50;
assign w254 = ~w50;
assign w255 = ~w51;
assign w256 = ~w51;
assign w257 = ~w51;
assign w258 = ~w52;
assign w259 = ~w52;
assign w260 = ~w52;
assign w261 = ~w53;
assign w262 = ~w54;
assign w263 = ~w55;
assign w264 = ~w55;
assign w265 = w53 | w56;
assign w266 = ~w56;
assign w267 = ~w57;
assign w268 = ~w57;
assign w269 = ~w59;
assign w270 = ~w59;
assign w271 = ~w60;
assign w272 = ~w61;
assign w273 = ~w62;
assign w274 = ~w62;
assign w275 = ~w63;
assign w276 = ~w63;
assign w277 = ~w64;
assign w278 = ~w64;
assign w279 = ~w65;
assign w280 = ~w65;
assign w281 = ~w66;
assign w282 = ~w66;
assign w283 = ~w67;
assign w284 = ~w67;
assign w285 = ~w68;
assign w286 = ~w68;
assign w287 = ~w69;
assign w288 = ~w69;
assign w289 = ~w70;
assign w290 = ~w70;
assign w291 = ~w71;
assign w292 = ~w71;
assign w293 = ~w72;
assign w294 = ~w72;
assign w295 = ~w73;
assign w296 = ~w73;
assign w297 = ~w74;
assign w298 = ~w74;
assign w299 = ~w75;
assign w300 = ~w75;
assign w301 = ~w76;
assign w302 = ~w76;
assign w303 = ~w77;
assign w304 = ~w77;
assign w305 = ~w78;
assign w306 = ~w78;
assign w307 = ~w79;
assign w308 = ~w79;
assign w309 = ~w84;
assign w310 = w80 & w86;
assign w311 = w80 ~^ w86;
assign w312 = ~w87;
assign w313 = w85 & w88;
assign w314 = w85 ~^ w88;
assign w315 = ~w89;
assign w316 = ~w89;
assign w317 = ~w90;
assign w318 = ~w90;
assign w319 = ~w90;
assign w320 = ~w91;
assign w321 = ~w91;
assign w322 = ~w91;
assign w323 = ~w92;
assign w324 = ~w93;
assign w325 = ~w94;
assign w326 = ~w94;
assign w327 = w92 | w95;
assign w328 = ~w95;
assign w329 = ~w96;
assign w330 = ~w96;
assign w331 = ~w98;
assign w332 = ~w98;
assign w333 = ~w99;
assign w334 = ~w100;
assign w335 = ~w101;
assign w336 = ~w101;
assign w337 = ~w102;
assign w338 = ~w102;
assign w339 = ~w103;
assign w340 = ~w103;
assign w341 = ~w104;
assign w342 = ~w104;
assign w343 = ~w105;
assign w344 = ~w105;
assign w345 = ~w106;
assign w346 = ~w106;
assign w347 = ~w107;
assign w348 = ~w107;
assign w349 = ~w108;
assign w350 = ~w108;
assign w351 = ~w109;
assign w352 = ~w109;
assign w353 = ~w114;
assign w354 = w110 & w116;
assign w355 = w110 ~^ w116;
assign w356 = ~w117;
assign w357 = w115 & w118;
assign w358 = w115 ~^ w118;
assign w359 = ~w119;
assign w360 = ~w119;
assign w361 = ~w120;
assign w362 = ~w120;
assign w363 = ~w120;
assign w364 = ~w121;
assign w365 = ~w121;
assign w366 = ~w121;
assign w367 = ~w122;
assign w368 = ~w123;
assign w369 = ~w124;
assign w370 = ~w124;
assign w371 = w122 | w125;
assign w372 = ~w125;
assign w373 = ~w126;
assign w374 = ~w126;
assign w375 = ~w128;
assign w376 = ~w128;
assign w377 = ~w133;
assign w378 = w129 & w135;
assign w379 = w129 ~^ w135;
assign w380 = ~w136;
assign w381 = w134 & w137;
assign w382 = w134 ~^ w137;
assign w383 = ~w138;
assign w384 = ~w138;
assign w385 = ~w139;
assign w386 = ~w139;
assign w387 = ~w139;
assign w388 = ~w140;
assign w389 = ~w140;
assign w390 = ~w140;
assign w391 = ~w141;
assign w392 = ~w142;
assign w393 = ~w143;
assign w394 = ~w143;
assign w395 = w141 | w144;
assign w396 = ~w144;
assign w397 = ~w145;
assign w398 = ~w145;
assign w399 = ~w147;
assign w400 = ~w147;
assign w401 = ~w148;
assign w402 = ~w149;
assign w403 = ~w153;
assign w404 = ~w154;
assign w405 = ~w155;
assign w406 = ~w155;
assign w407 = ~w156;
assign w408 = ~w156;
assign w409 = ~w157;
assign w410 = ~w157;
assign w411 = ~w158;
assign w412 = ~w158;
assign w413 = ~w159;
assign w414 = ~w159;
assign w415 = ~w160;
assign w416 = ~w160;
assign w417 = ~w161;
assign w418 = ~w161;
assign w419 = ~w162;
assign w420 = ~w162;
assign w421 = ~w163;
assign w422 = ~w163;
assign w423 = ~w168;
assign w424 = w164 & w170;
assign w425 = w164 ~^ w170;
assign w426 = ~w171;
assign w427 = w169 & w172;
assign w428 = w169 ~^ w172;
assign w429 = ~w173;
assign w430 = ~w173;
assign w431 = ~w174;
assign w432 = ~w174;
assign w433 = ~w174;
assign w434 = ~w175;
assign w435 = ~w175;
assign w436 = ~w175;
assign w437 = ~w176;
assign w438 = ~w177;
assign w439 = ~w178;
assign w440 = ~w178;
assign w441 = w176 | w179;
assign w442 = ~w179;
assign w443 = ~w180;
assign w444 = ~w180;
assign w445 = ~w182;
assign w446 = ~w182;
assign w447 = ~w183;
assign w448 = ~w183;
assign w449 = ~w184;
assign w450 = ~w184;
assign w451 = ~w185;
assign w452 = ~w186;
assign w453 = ~w186;
assign w454 = ~w187;
assign w455 = ~w187;
assign w456 = ~w188;
assign w457 = ~w188;
assign w458 = ~w189;
assign w459 = ~w189;
assign w460 = ~w190;
assign w461 = ~w191;
assign w462 = ~w192;
assign w463 = ~w192;
assign w464 = ~w193;
assign w465 = ~w194;
assign w466 = ~w194;
assign w467 = ~w195;
assign w468 = ~w195;
assign w469 = ~w196;
assign w470 = ~w197;
assign w471 = ~w197;
assign w472 = ~w198;
assign w473 = ~w199;
assign w474 = ~w199;
assign w475 = ~w200;
assign w476 = ~w201;
assign w477 = ~w202;
assign w478 = ~w202;
assign w479 = ~w203;
assign w480 = ~w204;
assign w481 = ~w206;
assign w482 = ~w206;
assign w483 = ~w207;
assign w484 = ~w209;
assign w485 = ~w209;
assign w486 = ~w210;
assign w487 = ~w210;
assign w488 = ~w211;
assign w489 = ~w212;
assign w490 = ~w212;
assign w491 = ~w213;
assign w492 = ~w213;
assign w493 = ~w214;
assign w494 = ~w215;
assign w495 = ~w215;
assign w496 = ~w216;
assign w497 = ~w216;
assign w498 = w205 ~^ w218;
assign w499 = ~w219;
assign w500 = ~w219;
assign w501 = ~w220;
assign w502 = w217 ~^ w222;
assign w503 = w217 ~| w222;
assign w504 = ~w223;
assign w505 = ~w223;
assign w506 = ~w224;
assign w507 = ~w224;
assign w508 = ~w225;
assign w509 = ~w225;
assign w510 = ~w226;
assign w511 = ~w226;
assign w512 = ~w227;
assign w513 = ~w227;
assign w514 = ~w228;
assign w515 = ~w228;
assign w516 = ~w229;
assign w517 = ~w230;
assign w518 = ~w230;
assign w519 = ~w231;
assign w520 = ~w231;
assign w521 = ~w232;
assign w522 = ~w232;
assign w523 = ~w233;
assign w524 = ~w233;
assign w525 = ~w234;
assign w526 = ~w235;
assign w527 = ~w236;
assign w528 = ~w236;
assign w529 = ~w237;
assign w530 = ~w238;
assign w531 = ~w238;
assign w532 = ~w239;
assign w533 = ~w239;
assign w534 = ~w240;
assign w535 = ~w241;
assign w536 = ~w241;
assign w537 = ~w242;
assign w538 = ~w243;
assign w539 = ~w243;
assign w540 = ~w244;
assign w541 = ~w245;
assign w542 = ~w246;
assign w543 = ~w246;
assign w544 = ~w247;
assign w545 = ~w248;
assign w546 = ~w250;
assign w547 = ~w250;
assign w548 = ~w251;
assign w549 = ~w253;
assign w550 = ~w253;
assign w551 = ~w254;
assign w552 = ~w254;
assign w553 = ~w255;
assign w554 = ~w256;
assign w555 = ~w256;
assign w556 = ~w257;
assign w557 = ~w257;
assign w558 = ~w258;
assign w559 = ~w259;
assign w560 = ~w259;
assign w561 = ~w260;
assign w562 = ~w260;
assign w563 = w249 ~^ w262;
assign w564 = ~w263;
assign w565 = ~w263;
assign w566 = ~w264;
assign w567 = w261 ~^ w266;
assign w568 = w261 ~| w266;
assign w569 = ~w267;
assign w570 = ~w267;
assign w571 = ~w268;
assign w572 = ~w268;
assign w573 = ~w269;
assign w574 = ~w269;
assign w575 = ~w270;
assign w576 = ~w270;
assign w577 = ~w271;
assign w578 = ~w271;
assign w579 = ~w272;
assign w580 = ~w272;
assign w581 = ~w273;
assign w582 = ~w274;
assign w583 = ~w274;
assign w584 = ~w275;
assign w585 = ~w275;
assign w586 = ~w276;
assign w587 = ~w276;
assign w588 = ~w277;
assign w589 = ~w277;
assign w590 = ~w278;
assign w591 = ~w279;
assign w592 = ~w280;
assign w593 = ~w280;
assign w594 = ~w281;
assign w595 = ~w282;
assign w596 = ~w282;
assign w597 = ~w283;
assign w598 = ~w283;
assign w599 = ~w284;
assign w600 = ~w285;
assign w601 = ~w285;
assign w602 = ~w286;
assign w603 = ~w287;
assign w604 = ~w287;
assign w605 = ~w288;
assign w606 = ~w289;
assign w607 = ~w290;
assign w608 = ~w290;
assign w609 = ~w291;
assign w610 = ~w292;
assign w611 = ~w292;
assign w612 = ~w293;
assign w613 = ~w293;
assign w614 = ~w294;
assign w615 = ~w294;
assign w616 = ~w295;
assign w617 = ~w295;
assign w618 = ~w296;
assign w619 = ~w297;
assign w620 = ~w298;
assign w621 = ~w298;
assign w622 = ~w299;
assign w623 = ~w300;
assign w624 = ~w300;
assign w625 = ~w301;
assign w626 = ~w301;
assign w627 = ~w302;
assign w628 = ~w303;
assign w629 = ~w303;
assign w630 = ~w304;
assign w631 = ~w305;
assign w632 = ~w305;
assign w633 = ~w306;
assign w634 = ~w307;
assign w635 = ~w308;
assign w636 = ~w308;
assign w637 = ~w309;
assign w638 = ~w310;
assign w639 = ~w312;
assign w640 = ~w312;
assign w641 = ~w313;
assign w642 = ~w315;
assign w643 = ~w315;
assign w644 = ~w316;
assign w645 = ~w316;
assign w646 = ~w317;
assign w647 = ~w318;
assign w648 = ~w318;
assign w649 = ~w319;
assign w650 = ~w319;
assign w651 = ~w320;
assign w652 = ~w321;
assign w653 = ~w321;
assign w654 = ~w322;
assign w655 = ~w322;
assign w656 = w311 ~^ w324;
assign w657 = ~w325;
assign w658 = ~w325;
assign w659 = ~w326;
assign w660 = w323 ~^ w328;
assign w661 = w323 ~| w328;
assign w662 = ~w329;
assign w663 = ~w329;
assign w664 = ~w330;
assign w665 = ~w330;
assign w666 = ~w331;
assign w667 = ~w331;
assign w668 = ~w332;
assign w669 = ~w332;
assign w670 = ~w333;
assign w671 = ~w333;
assign w672 = ~w334;
assign w673 = ~w334;
assign w674 = ~w335;
assign w675 = ~w336;
assign w676 = ~w336;
assign w677 = ~w337;
assign w678 = ~w337;
assign w679 = ~w338;
assign w680 = ~w338;
assign w681 = ~w339;
assign w682 = ~w339;
assign w683 = ~w340;
assign w684 = ~w341;
assign w685 = ~w342;
assign w686 = ~w342;
assign w687 = ~w343;
assign w688 = ~w344;
assign w689 = ~w344;
assign w690 = ~w345;
assign w691 = ~w345;
assign w692 = ~w346;
assign w693 = ~w347;
assign w694 = ~w347;
assign w695 = ~w348;
assign w696 = ~w349;
assign w697 = ~w349;
assign w698 = ~w350;
assign w699 = ~w351;
assign w700 = ~w352;
assign w701 = ~w352;
assign w702 = ~w353;
assign w703 = ~w354;
assign w704 = ~w356;
assign w705 = ~w356;
assign w706 = ~w357;
assign w707 = ~w359;
assign w708 = ~w359;
assign w709 = ~w360;
assign w710 = ~w360;
assign w711 = ~w361;
assign w712 = ~w362;
assign w713 = ~w362;
assign w714 = ~w363;
assign w715 = ~w363;
assign w716 = ~w364;
assign w717 = ~w365;
assign w718 = ~w365;
assign w719 = ~w366;
assign w720 = ~w366;
assign w721 = w355 ~^ w368;
assign w722 = ~w369;
assign w723 = ~w369;
assign w724 = ~w370;
assign w725 = w367 ~^ w372;
assign w726 = w367 ~| w372;
assign w727 = ~w373;
assign w728 = ~w373;
assign w729 = ~w374;
assign w730 = ~w374;
assign w731 = ~w375;
assign w732 = ~w375;
assign w733 = ~w376;
assign w734 = ~w376;
assign w735 = ~w377;
assign w736 = ~w378;
assign w737 = ~w380;
assign w738 = ~w380;
assign w739 = ~w381;
assign w740 = ~w383;
assign w741 = ~w383;
assign w742 = ~w384;
assign w743 = ~w384;
assign w744 = ~w385;
assign w745 = ~w386;
assign w746 = ~w386;
assign w747 = ~w387;
assign w748 = ~w387;
assign w749 = ~w388;
assign w750 = ~w389;
assign w751 = ~w389;
assign w752 = ~w390;
assign w753 = ~w390;
assign w754 = w379 ~^ w392;
assign w755 = ~w393;
assign w756 = ~w393;
assign w757 = ~w394;
assign w758 = w391 ~^ w396;
assign w759 = w391 ~| w396;
assign w760 = ~w397;
assign w761 = ~w397;
assign w762 = ~w398;
assign w763 = ~w398;
assign w764 = ~w399;
assign w765 = ~w399;
assign w766 = ~w400;
assign w767 = ~w400;
assign w768 = ~w401;
assign w769 = ~w401;
assign w770 = ~w402;
assign w771 = ~w402;
assign w772 = ~w403;
assign w773 = ~w403;
assign w774 = ~w404;
assign w775 = ~w404;
assign w776 = ~w405;
assign w777 = ~w406;
assign w778 = ~w406;
assign w779 = ~w407;
assign w780 = ~w407;
assign w781 = ~w408;
assign w782 = ~w408;
assign w783 = ~w409;
assign w784 = ~w409;
assign w785 = ~w410;
assign w786 = ~w411;
assign w787 = ~w412;
assign w788 = ~w412;
assign w789 = ~w413;
assign w790 = ~w414;
assign w791 = ~w414;
assign w792 = ~w415;
assign w793 = ~w415;
assign w794 = ~w416;
assign w795 = ~w417;
assign w796 = ~w417;
assign w797 = ~w418;
assign w798 = ~w419;
assign w799 = ~w419;
assign w800 = ~w420;
assign w801 = ~w421;
assign w802 = ~w422;
assign w803 = ~w422;
assign w804 = ~w423;
assign w805 = ~w424;
assign w806 = ~w426;
assign w807 = ~w426;
assign w808 = ~w427;
assign w809 = ~w429;
assign w810 = ~w429;
assign w811 = ~w430;
assign w812 = ~w430;
assign w813 = ~w431;
assign w814 = ~w432;
assign w815 = ~w432;
assign w816 = ~w433;
assign w817 = ~w433;
assign w818 = ~w434;
assign w819 = ~w435;
assign w820 = ~w435;
assign w821 = ~w436;
assign w822 = ~w436;
assign w823 = w425 ~^ w438;
assign w824 = ~w439;
assign w825 = ~w439;
assign w826 = ~w440;
assign w827 = w437 ~^ w442;
assign w828 = w437 ~| w442;
assign w829 = ~w443;
assign w830 = ~w443;
assign w831 = ~w444;
assign w832 = ~w444;
assign w833 = ~w445;
assign w834 = ~w445;
assign w835 = ~w446;
assign w836 = ~w446;
assign w837 = ~w447;
assign w838 = ~w447;
assign w839 = ~w448;
assign w840 = ~w448;
assign w841 = ~w449;
assign w842 = ~w449;
assign w843 = ~w450;
assign w844 = ~w450;
assign w845 = ~w451;
assign w846 = w15 | w460;
assign w847 = w25 | w468;
assign w848 = ~w479;
assign w849 = ~w481;
assign w850 = ~w482;
assign w851 = w464 | w484;
assign w852 = w462 | w484;
assign w853 = w469 | w485;
assign w854 = w458 | w486;
assign w855 = w476 | w486;
assign w856 = w470 | w487;
assign w857 = w454 | w487;
assign w858 = w467 | w488;
assign w859 = w478 | w488;
assign w860 = w459 | w489;
assign w861 = w6 | w489;
assign w862 = w470 | w490;
assign w863 = w453 | w490;
assign w864 = w456 | w491;
assign w865 = w474 | w491;
assign w866 = w462 | w492;
assign w867 = w466 | w493;
assign w868 = w477 | w493;
assign w869 = w7 | w494;
assign w870 = w9 | w494;
assign w871 = w4 | w495;
assign w872 = w472 | w495;
assign w873 = w455 | w496;
assign w874 = w461 | w496;
assign w875 = w457 | w499;
assign w876 = w10 | w499;
assign w877 = w465 | w500;
assign w878 = w460 | w500;
assign w879 = w473 | w501;
assign w880 = w471 | w501;
assign w881 = w469 | w504;
assign w882 = w474 | w504;
assign w883 = w465 | w505;
assign w884 = w453 | w505;
assign w885 = w463 | w506;
assign w886 = w457 | w506;
assign w887 = w477 | w507;
assign w888 = w471 | w507;
assign w889 = w468 | w508;
assign w890 = w464 | w508;
assign w891 = w473 | w509;
assign w892 = w455 | w509;
assign w893 = w8 | w510;
assign w894 = w459 | w510;
assign w895 = w5 | w511;
assign w896 = w452 | w511;
assign w897 = ~w512;
assign w898 = ~w512;
assign w899 = ~w513;
assign w900 = ~w513;
assign w901 = ~w514;
assign w902 = ~w514;
assign w903 = ~w515;
assign w904 = ~w515;
assign w905 = ~w516;
assign w906 = w45 | w525;
assign w907 = w55 | w533;
assign w908 = ~w544;
assign w909 = ~w546;
assign w910 = ~w547;
assign w911 = w529 | w549;
assign w912 = w527 | w549;
assign w913 = w534 | w550;
assign w914 = w523 | w551;
assign w915 = w541 | w551;
assign w916 = w535 | w552;
assign w917 = w519 | w552;
assign w918 = w532 | w553;
assign w919 = w543 | w553;
assign w920 = w524 | w554;
assign w921 = w36 | w554;
assign w922 = w535 | w555;
assign w923 = w518 | w555;
assign w924 = w521 | w556;
assign w925 = w539 | w556;
assign w926 = w527 | w557;
assign w927 = w531 | w558;
assign w928 = w542 | w558;
assign w929 = w37 | w559;
assign w930 = w39 | w559;
assign w931 = w34 | w560;
assign w932 = w537 | w560;
assign w933 = w520 | w561;
assign w934 = w526 | w561;
assign w935 = w522 | w564;
assign w936 = w40 | w564;
assign w937 = w530 | w565;
assign w938 = w525 | w565;
assign w939 = w538 | w566;
assign w940 = w536 | w566;
assign w941 = w534 | w569;
assign w942 = w539 | w569;
assign w943 = w530 | w570;
assign w944 = w518 | w570;
assign w945 = w528 | w571;
assign w946 = w522 | w571;
assign w947 = w542 | w572;
assign w948 = w536 | w572;
assign w949 = w533 | w573;
assign w950 = w529 | w573;
assign w951 = w538 | w574;
assign w952 = w520 | w574;
assign w953 = w38 | w575;
assign w954 = w524 | w575;
assign w955 = w35 | w576;
assign w956 = w517 | w576;
assign w957 = ~w577;
assign w958 = ~w577;
assign w959 = ~w578;
assign w960 = ~w578;
assign w961 = ~w579;
assign w962 = ~w579;
assign w963 = ~w580;
assign w964 = ~w580;
assign w965 = ~w581;
assign w966 = w133 | w590;
assign w967 = w143 | w598;
assign w968 = ~w609;
assign w969 = w84 | w618;
assign w970 = w94 | w626;
assign w971 = ~w637;
assign w972 = ~w639;
assign w973 = ~w640;
assign w974 = w622 | w642;
assign w975 = w620 | w642;
assign w976 = w627 | w643;
assign w977 = w616 | w644;
assign w978 = w634 | w644;
assign w979 = w628 | w645;
assign w980 = w612 | w645;
assign w981 = w625 | w646;
assign w982 = w636 | w646;
assign w983 = w617 | w647;
assign w984 = w75 | w647;
assign w985 = w628 | w648;
assign w986 = w611 | w648;
assign w987 = w614 | w649;
assign w988 = w632 | w649;
assign w989 = w620 | w650;
assign w990 = w624 | w651;
assign w991 = w635 | w651;
assign w992 = w76 | w652;
assign w993 = w78 | w652;
assign w994 = w73 | w653;
assign w995 = w630 | w653;
assign w996 = w613 | w654;
assign w997 = w619 | w654;
assign w998 = w615 | w657;
assign w999 = w79 | w657;
assign w1000 = w623 | w658;
assign w1001 = w618 | w658;
assign w1002 = w631 | w659;
assign w1003 = w629 | w659;
assign w1004 = w627 | w662;
assign w1005 = w632 | w662;
assign w1006 = w623 | w663;
assign w1007 = w611 | w663;
assign w1008 = w621 | w664;
assign w1009 = w615 | w664;
assign w1010 = w635 | w665;
assign w1011 = w629 | w665;
assign w1012 = w626 | w666;
assign w1013 = w622 | w666;
assign w1014 = w631 | w667;
assign w1015 = w613 | w667;
assign w1016 = w77 | w668;
assign w1017 = w617 | w668;
assign w1018 = w74 | w669;
assign w1019 = w610 | w669;
assign w1020 = ~w670;
assign w1021 = ~w670;
assign w1022 = ~w671;
assign w1023 = ~w671;
assign w1024 = ~w672;
assign w1025 = ~w672;
assign w1026 = ~w673;
assign w1027 = ~w673;
assign w1028 = ~w674;
assign w1029 = w114 | w683;
assign w1030 = w124 | w691;
assign w1031 = ~w702;
assign w1032 = ~w704;
assign w1033 = ~w705;
assign w1034 = w687 | w707;
assign w1035 = w685 | w707;
assign w1036 = w692 | w708;
assign w1037 = w681 | w709;
assign w1038 = w699 | w709;
assign w1039 = w693 | w710;
assign w1040 = w677 | w710;
assign w1041 = w690 | w711;
assign w1042 = w701 | w711;
assign w1043 = w682 | w712;
assign w1044 = w105 | w712;
assign w1045 = w693 | w713;
assign w1046 = w676 | w713;
assign w1047 = w679 | w714;
assign w1048 = w697 | w714;
assign w1049 = w685 | w715;
assign w1050 = w689 | w716;
assign w1051 = w700 | w716;
assign w1052 = w106 | w717;
assign w1053 = w108 | w717;
assign w1054 = w103 | w718;
assign w1055 = w695 | w718;
assign w1056 = w678 | w719;
assign w1057 = w684 | w719;
assign w1058 = w680 | w722;
assign w1059 = w109 | w722;
assign w1060 = w688 | w723;
assign w1061 = w683 | w723;
assign w1062 = w696 | w724;
assign w1063 = w694 | w724;
assign w1064 = w692 | w727;
assign w1065 = w697 | w727;
assign w1066 = w688 | w728;
assign w1067 = w676 | w728;
assign w1068 = w686 | w729;
assign w1069 = w680 | w729;
assign w1070 = w700 | w730;
assign w1071 = w694 | w730;
assign w1072 = w691 | w731;
assign w1073 = w687 | w731;
assign w1074 = w696 | w732;
assign w1075 = w678 | w732;
assign w1076 = w107 | w733;
assign w1077 = w682 | w733;
assign w1078 = w104 | w734;
assign w1079 = w675 | w734;
assign w1080 = ~w735;
assign w1081 = ~w737;
assign w1082 = ~w738;
assign w1083 = w594 | w740;
assign w1084 = w592 | w740;
assign w1085 = w599 | w741;
assign w1086 = w588 | w742;
assign w1087 = w606 | w742;
assign w1088 = w600 | w743;
assign w1089 = w584 | w743;
assign w1090 = w597 | w744;
assign w1091 = w608 | w744;
assign w1092 = w589 | w745;
assign w1093 = w66 | w745;
assign w1094 = w600 | w746;
assign w1095 = w583 | w746;
assign w1096 = w586 | w747;
assign w1097 = w604 | w747;
assign w1098 = w592 | w748;
assign w1099 = w596 | w749;
assign w1100 = w607 | w749;
assign w1101 = w67 | w750;
assign w1102 = w69 | w750;
assign w1103 = w64 | w751;
assign w1104 = w602 | w751;
assign w1105 = w585 | w752;
assign w1106 = w591 | w752;
assign w1107 = w587 | w755;
assign w1108 = w70 | w755;
assign w1109 = w595 | w756;
assign w1110 = w590 | w756;
assign w1111 = w603 | w757;
assign w1112 = w601 | w757;
assign w1113 = w599 | w760;
assign w1114 = w604 | w760;
assign w1115 = w595 | w761;
assign w1116 = w583 | w761;
assign w1117 = w593 | w762;
assign w1118 = w587 | w762;
assign w1119 = w607 | w763;
assign w1120 = w601 | w763;
assign w1121 = w598 | w764;
assign w1122 = w594 | w764;
assign w1123 = w603 | w765;
assign w1124 = w585 | w765;
assign w1125 = w68 | w766;
assign w1126 = w589 | w766;
assign w1127 = w65 | w767;
assign w1128 = w582 | w767;
assign w1129 = ~w768;
assign w1130 = ~w768;
assign w1131 = ~w769;
assign w1132 = ~w769;
assign w1133 = ~w770;
assign w1134 = ~w770;
assign w1135 = ~w771;
assign w1136 = ~w771;
assign w1137 = ~w772;
assign w1138 = ~w772;
assign w1139 = ~w773;
assign w1140 = ~w773;
assign w1141 = ~w774;
assign w1142 = ~w774;
assign w1143 = ~w775;
assign w1144 = ~w775;
assign w1145 = ~w776;
assign w1146 = w168 | w785;
assign w1147 = w178 | w793;
assign w1148 = ~w804;
assign w1149 = ~w806;
assign w1150 = ~w807;
assign w1151 = w789 | w809;
assign w1152 = w787 | w809;
assign w1153 = w794 | w810;
assign w1154 = w783 | w811;
assign w1155 = w801 | w811;
assign w1156 = w795 | w812;
assign w1157 = w779 | w812;
assign w1158 = w792 | w813;
assign w1159 = w803 | w813;
assign w1160 = w784 | w814;
assign w1161 = w159 | w814;
assign w1162 = w795 | w815;
assign w1163 = w778 | w815;
assign w1164 = w781 | w816;
assign w1165 = w799 | w816;
assign w1166 = w787 | w817;
assign w1167 = w791 | w818;
assign w1168 = w802 | w818;
assign w1169 = w160 | w819;
assign w1170 = w162 | w819;
assign w1171 = w157 | w820;
assign w1172 = w797 | w820;
assign w1173 = w780 | w821;
assign w1174 = w786 | w821;
assign w1175 = w782 | w824;
assign w1176 = w163 | w824;
assign w1177 = w790 | w825;
assign w1178 = w785 | w825;
assign w1179 = w798 | w826;
assign w1180 = w796 | w826;
assign w1181 = w794 | w829;
assign w1182 = w799 | w829;
assign w1183 = w790 | w830;
assign w1184 = w778 | w830;
assign w1185 = w788 | w831;
assign w1186 = w782 | w831;
assign w1187 = w802 | w832;
assign w1188 = w796 | w832;
assign w1189 = w793 | w833;
assign w1190 = w789 | w833;
assign w1191 = w798 | w834;
assign w1192 = w780 | w834;
assign w1193 = w161 | w835;
assign w1194 = w784 | w835;
assign w1195 = w158 | w836;
assign w1196 = w777 | w836;
assign w1197 = ~w837;
assign w1198 = ~w837;
assign w1199 = ~w838;
assign w1200 = ~w838;
assign w1201 = ~w839;
assign w1202 = ~w839;
assign w1203 = ~w840;
assign w1204 = ~w840;
assign w1205 = ~w841;
assign w1206 = ~w841;
assign w1207 = ~w842;
assign w1208 = ~w842;
assign w1209 = ~w843;
assign w1210 = ~w843;
assign w1211 = ~w844;
assign w1212 = ~w844;
assign w1213 = ~w845;
assign w1214 = ~w845;
assign w1215 = ~w848;
assign w1216 = ~w848;
assign w1217 = ~w849;
assign w1218 = ~w849;
assign w1219 = ~w850;
assign w1220 = ~w850;
assign w1221 = w857 ~^ w863;
assign w1222 = w857 & w863;
assign w1223 = w857 ~| w863;
assign w1224 = w855 ~^ w865;
assign w1225 = w847 | w865;
assign w1226 = w847 & w865;
assign w1227 = w859 ~^ w870;
assign w1228 = w866 ~^ w871;
assign w1229 = w866 | w871;
assign w1230 = w866 & w871;
assign w1231 = w860 ~^ w873;
assign w1232 = w860 & w873;
assign w1233 = w860 | w873;
assign w1234 = w869 ~^ w877;
assign w1235 = w869 & w877;
assign w1236 = w869 | w877;
assign w1237 = w853 ~^ w878;
assign w1238 = w868 ~^ w879;
assign w1239 = w870 & w881;
assign w1240 = w870 | w881;
assign w1241 = w876 ~^ w882;
assign w1242 = w872 ~^ w883;
assign w1243 = w875 ~^ w884;
assign w1244 = w875 & w884;
assign w1245 = w875 | w884;
assign w1246 = w878 | w886;
assign w1247 = w878 & w886;
assign w1248 = w879 | w889;
assign w1249 = w879 & w889;
assign w1250 = w880 ~^ w890;
assign w1251 = w880 | w890;
assign w1252 = w880 & w890;
assign w1253 = w887 ~^ w891;
assign w1254 = w887 & w891;
assign w1255 = w887 ~| w891;
assign w1256 = w867 ~^ w892;
assign w1257 = w867 | w892;
assign w1258 = w867 & w892;
assign w1259 = w882 & w893;
assign w1260 = w882 | w893;
assign w1261 = w885 ~^ w894;
assign w1262 = w885 & w894;
assign w1263 = w885 | w894;
assign w1264 = w883 | w895;
assign w1265 = w883 & w895;
assign w1266 = w861 ~^ w896;
assign w1267 = w874 & w896;
assign w1268 = w874 | w896;
assign w1269 = ~w897;
assign w1270 = ~w897;
assign w1271 = ~w898;
assign w1272 = ~w898;
assign w1273 = ~w899;
assign w1274 = ~w899;
assign w1275 = ~w900;
assign w1276 = ~w900;
assign w1277 = ~w901;
assign w1278 = ~w901;
assign w1279 = ~w902;
assign w1280 = ~w902;
assign w1281 = ~w903;
assign w1282 = ~w903;
assign w1283 = ~w904;
assign w1284 = ~w904;
assign w1285 = ~w905;
assign w1286 = ~w905;
assign w1287 = ~w908;
assign w1288 = ~w908;
assign w1289 = ~w909;
assign w1290 = ~w909;
assign w1291 = ~w910;
assign w1292 = ~w910;
assign w1293 = w917 ~^ w923;
assign w1294 = w917 & w923;
assign w1295 = w917 ~| w923;
assign w1296 = w915 ~^ w925;
assign w1297 = w907 | w925;
assign w1298 = w907 & w925;
assign w1299 = w919 ~^ w930;
assign w1300 = w926 ~^ w931;
assign w1301 = w926 | w931;
assign w1302 = w926 & w931;
assign w1303 = w920 ~^ w933;
assign w1304 = w920 & w933;
assign w1305 = w920 | w933;
assign w1306 = w929 ~^ w937;
assign w1307 = w929 & w937;
assign w1308 = w929 | w937;
assign w1309 = w913 ~^ w938;
assign w1310 = w928 ~^ w939;
assign w1311 = w930 & w941;
assign w1312 = w930 | w941;
assign w1313 = w936 ~^ w942;
assign w1314 = w932 ~^ w943;
assign w1315 = w935 ~^ w944;
assign w1316 = w935 & w944;
assign w1317 = w935 | w944;
assign w1318 = w938 | w946;
assign w1319 = w938 & w946;
assign w1320 = w939 | w949;
assign w1321 = w939 & w949;
assign w1322 = w940 ~^ w950;
assign w1323 = w940 | w950;
assign w1324 = w940 & w950;
assign w1325 = w947 ~^ w951;
assign w1326 = w947 & w951;
assign w1327 = w947 ~| w951;
assign w1328 = w927 ~^ w952;
assign w1329 = w927 | w952;
assign w1330 = w927 & w952;
assign w1331 = w942 & w953;
assign w1332 = w942 | w953;
assign w1333 = w945 ~^ w954;
assign w1334 = w945 & w954;
assign w1335 = w945 | w954;
assign w1336 = w943 | w955;
assign w1337 = w943 & w955;
assign w1338 = w921 ~^ w956;
assign w1339 = w934 & w956;
assign w1340 = w934 | w956;
assign w1341 = ~w957;
assign w1342 = ~w957;
assign w1343 = ~w958;
assign w1344 = ~w958;
assign w1345 = ~w959;
assign w1346 = ~w959;
assign w1347 = ~w960;
assign w1348 = ~w960;
assign w1349 = ~w961;
assign w1350 = ~w961;
assign w1351 = ~w962;
assign w1352 = ~w962;
assign w1353 = ~w963;
assign w1354 = ~w963;
assign w1355 = ~w964;
assign w1356 = ~w964;
assign w1357 = ~w965;
assign w1358 = ~w965;
assign w1359 = ~w968;
assign w1360 = ~w968;
assign w1361 = ~w971;
assign w1362 = ~w971;
assign w1363 = ~w972;
assign w1364 = ~w972;
assign w1365 = ~w973;
assign w1366 = ~w973;
assign w1367 = w980 ~^ w986;
assign w1368 = w980 & w986;
assign w1369 = w980 ~| w986;
assign w1370 = w978 ~^ w988;
assign w1371 = w970 | w988;
assign w1372 = w970 & w988;
assign w1373 = w982 ~^ w993;
assign w1374 = w989 ~^ w994;
assign w1375 = w989 | w994;
assign w1376 = w989 & w994;
assign w1377 = w983 ~^ w996;
assign w1378 = w983 & w996;
assign w1379 = w983 | w996;
assign w1380 = w992 ~^ w1000;
assign w1381 = w992 & w1000;
assign w1382 = w992 | w1000;
assign w1383 = w976 ~^ w1001;
assign w1384 = w991 ~^ w1002;
assign w1385 = w993 & w1004;
assign w1386 = w993 | w1004;
assign w1387 = w999 ~^ w1005;
assign w1388 = w995 ~^ w1006;
assign w1389 = w998 ~^ w1007;
assign w1390 = w998 & w1007;
assign w1391 = w998 | w1007;
assign w1392 = w1001 | w1009;
assign w1393 = w1001 & w1009;
assign w1394 = w1002 | w1012;
assign w1395 = w1002 & w1012;
assign w1396 = w1003 ~^ w1013;
assign w1397 = w1003 | w1013;
assign w1398 = w1003 & w1013;
assign w1399 = w1010 ~^ w1014;
assign w1400 = w1010 & w1014;
assign w1401 = w1010 ~| w1014;
assign w1402 = w990 ~^ w1015;
assign w1403 = w990 | w1015;
assign w1404 = w990 & w1015;
assign w1405 = w1005 & w1016;
assign w1406 = w1005 | w1016;
assign w1407 = w1008 ~^ w1017;
assign w1408 = w1008 & w1017;
assign w1409 = w1008 | w1017;
assign w1410 = w1006 | w1018;
assign w1411 = w1006 & w1018;
assign w1412 = w984 ~^ w1019;
assign w1413 = w997 & w1019;
assign w1414 = w997 | w1019;
assign w1415 = ~w1020;
assign w1416 = ~w1020;
assign w1417 = ~w1021;
assign w1418 = ~w1021;
assign w1419 = ~w1022;
assign w1420 = ~w1022;
assign w1421 = ~w1023;
assign w1422 = ~w1023;
assign w1423 = ~w1024;
assign w1424 = ~w1024;
assign w1425 = ~w1025;
assign w1426 = ~w1025;
assign w1427 = ~w1026;
assign w1428 = ~w1026;
assign w1429 = ~w1027;
assign w1430 = ~w1027;
assign w1431 = ~w1028;
assign w1432 = ~w1028;
assign w1433 = ~w1031;
assign w1434 = ~w1031;
assign w1435 = ~w1032;
assign w1436 = ~w1032;
assign w1437 = ~w1033;
assign w1438 = ~w1033;
assign w1439 = w1040 ~^ w1046;
assign w1440 = w1040 & w1046;
assign w1441 = w1040 ~| w1046;
assign w1442 = w1038 ~^ w1048;
assign w1443 = w1030 | w1048;
assign w1444 = w1030 & w1048;
assign w1445 = w1042 ~^ w1053;
assign w1446 = w1049 ~^ w1054;
assign w1447 = w1049 | w1054;
assign w1448 = w1049 & w1054;
assign w1449 = w1043 ~^ w1056;
assign w1450 = w1043 & w1056;
assign w1451 = w1043 | w1056;
assign w1452 = w1052 ~^ w1060;
assign w1453 = w1052 & w1060;
assign w1454 = w1052 | w1060;
assign w1455 = w1036 ~^ w1061;
assign w1456 = w1051 ~^ w1062;
assign w1457 = w1053 & w1064;
assign w1458 = w1053 | w1064;
assign w1459 = w1059 ~^ w1065;
assign w1460 = w1055 ~^ w1066;
assign w1461 = w1058 ~^ w1067;
assign w1462 = w1058 & w1067;
assign w1463 = w1058 | w1067;
assign w1464 = w1061 | w1069;
assign w1465 = w1061 & w1069;
assign w1466 = w1062 | w1072;
assign w1467 = w1062 & w1072;
assign w1468 = w1063 ~^ w1073;
assign w1469 = w1063 | w1073;
assign w1470 = w1063 & w1073;
assign w1471 = w1070 ~^ w1074;
assign w1472 = w1070 & w1074;
assign w1473 = w1070 ~| w1074;
assign w1474 = w1050 ~^ w1075;
assign w1475 = w1050 | w1075;
assign w1476 = w1050 & w1075;
assign w1477 = w1065 & w1076;
assign w1478 = w1065 | w1076;
assign w1479 = w1068 ~^ w1077;
assign w1480 = w1068 & w1077;
assign w1481 = w1068 | w1077;
assign w1482 = w1066 | w1078;
assign w1483 = w1066 & w1078;
assign w1484 = w1044 ~^ w1079;
assign w1485 = w1057 & w1079;
assign w1486 = w1057 | w1079;
assign w1487 = ~w1080;
assign w1488 = ~w1080;
assign w1489 = ~w1081;
assign w1490 = ~w1081;
assign w1491 = ~w1082;
assign w1492 = ~w1082;
assign w1493 = w1089 ~^ w1095;
assign w1494 = w1089 & w1095;
assign w1495 = w1089 ~| w1095;
assign w1496 = w1087 ~^ w1097;
assign w1497 = w967 | w1097;
assign w1498 = w967 & w1097;
assign w1499 = w1091 ~^ w1102;
assign w1500 = w1098 ~^ w1103;
assign w1501 = w1098 | w1103;
assign w1502 = w1098 & w1103;
assign w1503 = w1092 ~^ w1105;
assign w1504 = w1092 & w1105;
assign w1505 = w1092 | w1105;
assign w1506 = w1101 ~^ w1109;
assign w1507 = w1101 & w1109;
assign w1508 = w1101 | w1109;
assign w1509 = w1085 ~^ w1110;
assign w1510 = w1100 ~^ w1111;
assign w1511 = w1102 & w1113;
assign w1512 = w1102 | w1113;
assign w1513 = w1108 ~^ w1114;
assign w1514 = w1104 ~^ w1115;
assign w1515 = w1107 ~^ w1116;
assign w1516 = w1107 & w1116;
assign w1517 = w1107 | w1116;
assign w1518 = w1110 | w1118;
assign w1519 = w1110 & w1118;
assign w1520 = w1111 | w1121;
assign w1521 = w1111 & w1121;
assign w1522 = w1112 ~^ w1122;
assign w1523 = w1112 | w1122;
assign w1524 = w1112 & w1122;
assign w1525 = w1119 ~^ w1123;
assign w1526 = w1119 & w1123;
assign w1527 = w1119 ~| w1123;
assign w1528 = w1099 ~^ w1124;
assign w1529 = w1099 | w1124;
assign w1530 = w1099 & w1124;
assign w1531 = w1114 & w1125;
assign w1532 = w1114 | w1125;
assign w1533 = w1117 ~^ w1126;
assign w1534 = w1117 & w1126;
assign w1535 = w1117 | w1126;
assign w1536 = w1115 | w1127;
assign w1537 = w1115 & w1127;
assign w1538 = w1093 ~^ w1128;
assign w1539 = w1106 & w1128;
assign w1540 = w1106 | w1128;
assign w1541 = ~w1129;
assign w1542 = ~w1129;
assign w1543 = ~w1130;
assign w1544 = ~w1130;
assign w1545 = ~w1131;
assign w1546 = ~w1131;
assign w1547 = ~w1132;
assign w1548 = ~w1132;
assign w1549 = ~w1133;
assign w1550 = ~w1133;
assign w1551 = ~w1134;
assign w1552 = ~w1134;
assign w1553 = ~w1135;
assign w1554 = ~w1135;
assign w1555 = ~w1136;
assign w1556 = ~w1136;
assign w1557 = ~w1137;
assign w1558 = ~w1137;
assign w1559 = ~w1138;
assign w1560 = ~w1138;
assign w1561 = ~w1139;
assign w1562 = ~w1139;
assign w1563 = ~w1140;
assign w1564 = ~w1140;
assign w1565 = ~w1141;
assign w1566 = ~w1141;
assign w1567 = ~w1142;
assign w1568 = ~w1142;
assign w1569 = ~w1143;
assign w1570 = ~w1143;
assign w1571 = ~w1144;
assign w1572 = ~w1144;
assign w1573 = ~w1145;
assign w1574 = ~w1145;
assign w1575 = ~w1148;
assign w1576 = ~w1148;
assign w1577 = ~w1149;
assign w1578 = ~w1149;
assign w1579 = ~w1150;
assign w1580 = ~w1150;
assign w1581 = w1157 ~^ w1163;
assign w1582 = w1157 & w1163;
assign w1583 = w1157 ~| w1163;
assign w1584 = w1155 ~^ w1165;
assign w1585 = w1147 | w1165;
assign w1586 = w1147 & w1165;
assign w1587 = w1159 ~^ w1170;
assign w1588 = w1166 ~^ w1171;
assign w1589 = w1166 | w1171;
assign w1590 = w1166 & w1171;
assign w1591 = w1160 ~^ w1173;
assign w1592 = w1160 & w1173;
assign w1593 = w1160 | w1173;
assign w1594 = w1169 ~^ w1177;
assign w1595 = w1169 & w1177;
assign w1596 = w1169 | w1177;
assign w1597 = w1153 ~^ w1178;
assign w1598 = w1168 ~^ w1179;
assign w1599 = w1170 & w1181;
assign w1600 = w1170 | w1181;
assign w1601 = w1176 ~^ w1182;
assign w1602 = w1172 ~^ w1183;
assign w1603 = w1175 ~^ w1184;
assign w1604 = w1175 & w1184;
assign w1605 = w1175 | w1184;
assign w1606 = w1178 | w1186;
assign w1607 = w1178 & w1186;
assign w1608 = w1179 | w1189;
assign w1609 = w1179 & w1189;
assign w1610 = w1180 ~^ w1190;
assign w1611 = w1180 | w1190;
assign w1612 = w1180 & w1190;
assign w1613 = w1187 ~^ w1191;
assign w1614 = w1187 & w1191;
assign w1615 = w1187 ~| w1191;
assign w1616 = w1167 ~^ w1192;
assign w1617 = w1167 | w1192;
assign w1618 = w1167 & w1192;
assign w1619 = w1182 & w1193;
assign w1620 = w1182 | w1193;
assign w1621 = w1185 ~^ w1194;
assign w1622 = w1185 & w1194;
assign w1623 = w1185 | w1194;
assign w1624 = w1183 | w1195;
assign w1625 = w1183 & w1195;
assign w1626 = w1161 ~^ w1196;
assign w1627 = w1174 & w1196;
assign w1628 = w1174 | w1196;
assign w1629 = ~w1197;
assign w1630 = w28 & w1202;
assign w1631 = ~w1205;
assign w1632 = w15 ~| w1213;
assign w1633 = w497 | w1214;
assign w1634 = w485 | w1214;
assign w1635 = w454 ~| w1215;
assign w1636 = w476 | w1216;
assign w1637 = w475 | w1216;
assign w1638 = w452 ~| w1217;
assign w1639 = w475 | w1217;
assign w1640 = w472 | w1218;
assign w1641 = w461 | w1218;
assign w1642 = w456 ~| w1219;
assign w1643 = w458 | w1220;
assign w1644 = w467 | w1220;
assign w1645 = w847 ~^ w1224;
assign w1646 = w855 | w1226;
assign w1647 = w881 ~^ w1227;
assign w1648 = w851 ~^ w1228;
assign w1649 = w851 | w1230;
assign w1650 = w852 ~^ w1231;
assign w1651 = w852 | w1232;
assign w1652 = w862 ~^ w1234;
assign w1653 = w862 | w1235;
assign w1654 = w886 ~^ w1237;
assign w1655 = w889 ~^ w1238;
assign w1656 = w859 | w1239;
assign w1657 = w893 ~^ w1241;
assign w1658 = w895 ~^ w1242;
assign w1659 = w204 ~^ w1243;
assign w1660 = w480 | w1244;
assign w1661 = w853 | w1247;
assign w1662 = w868 | w1249;
assign w1663 = w856 ~^ w1256;
assign w1664 = w856 | w1258;
assign w1665 = w876 | w1259;
assign w1666 = w208 ~^ w1261;
assign w1667 = w208 | w1262;
assign w1668 = w872 | w1265;
assign w1669 = w874 ~^ w1266;
assign w1670 = w861 | w1267;
assign w1671 = ~w1269;
assign w1672 = w58 & w1274;
assign w1673 = ~w1277;
assign w1674 = w45 ~| w1285;
assign w1675 = w562 | w1286;
assign w1676 = w550 | w1286;
assign w1677 = w519 ~| w1287;
assign w1678 = w541 | w1288;
assign w1679 = w540 | w1288;
assign w1680 = w517 ~| w1289;
assign w1681 = w540 | w1289;
assign w1682 = w537 | w1290;
assign w1683 = w526 | w1290;
assign w1684 = w521 ~| w1291;
assign w1685 = w523 | w1292;
assign w1686 = w532 | w1292;
assign w1687 = w907 ~^ w1296;
assign w1688 = w915 | w1298;
assign w1689 = w941 ~^ w1299;
assign w1690 = w911 ~^ w1300;
assign w1691 = w911 | w1302;
assign w1692 = w912 ~^ w1303;
assign w1693 = w912 | w1304;
assign w1694 = w922 ~^ w1306;
assign w1695 = w922 | w1307;
assign w1696 = w946 ~^ w1309;
assign w1697 = w949 ~^ w1310;
assign w1698 = w919 | w1311;
assign w1699 = w953 ~^ w1313;
assign w1700 = w955 ~^ w1314;
assign w1701 = w248 ~^ w1315;
assign w1702 = w545 | w1316;
assign w1703 = w913 | w1319;
assign w1704 = w928 | w1321;
assign w1705 = w916 ~^ w1328;
assign w1706 = w916 | w1330;
assign w1707 = w936 | w1331;
assign w1708 = w252 ~^ w1333;
assign w1709 = w252 | w1334;
assign w1710 = w932 | w1337;
assign w1711 = w934 ~^ w1338;
assign w1712 = w921 | w1339;
assign w1713 = ~w1341;
assign w1714 = w97 & w1346;
assign w1715 = ~w1349;
assign w1716 = w133 ~| w1357;
assign w1717 = w753 | w1358;
assign w1718 = w741 | w1358;
assign w1719 = w84 ~| w1359;
assign w1720 = w655 | w1360;
assign w1721 = w643 | w1360;
assign w1722 = w612 ~| w1361;
assign w1723 = w634 | w1362;
assign w1724 = w633 | w1362;
assign w1725 = w610 ~| w1363;
assign w1726 = w633 | w1363;
assign w1727 = w630 | w1364;
assign w1728 = w619 | w1364;
assign w1729 = w614 ~| w1365;
assign w1730 = w616 | w1366;
assign w1731 = w625 | w1366;
assign w1732 = w970 ~^ w1370;
assign w1733 = w978 | w1372;
assign w1734 = w1004 ~^ w1373;
assign w1735 = w974 ~^ w1374;
assign w1736 = w974 | w1376;
assign w1737 = w975 ~^ w1377;
assign w1738 = w975 | w1378;
assign w1739 = w985 ~^ w1380;
assign w1740 = w985 | w1381;
assign w1741 = w1009 ~^ w1383;
assign w1742 = w1012 ~^ w1384;
assign w1743 = w982 | w1385;
assign w1744 = w1016 ~^ w1387;
assign w1745 = w1018 ~^ w1388;
assign w1746 = w310 ~^ w1389;
assign w1747 = w638 | w1390;
assign w1748 = w976 | w1393;
assign w1749 = w991 | w1395;
assign w1750 = w979 ~^ w1402;
assign w1751 = w979 | w1404;
assign w1752 = w999 | w1405;
assign w1753 = w314 ~^ w1407;
assign w1754 = w314 | w1408;
assign w1755 = w995 | w1411;
assign w1756 = w997 ~^ w1412;
assign w1757 = w984 | w1413;
assign w1758 = ~w1415;
assign w1759 = w127 & w1420;
assign w1760 = ~w1423;
assign w1761 = w114 ~| w1431;
assign w1762 = w720 | w1432;
assign w1763 = w708 | w1432;
assign w1764 = w677 ~| w1433;
assign w1765 = w699 | w1434;
assign w1766 = w698 | w1434;
assign w1767 = w675 ~| w1435;
assign w1768 = w698 | w1435;
assign w1769 = w695 | w1436;
assign w1770 = w684 | w1436;
assign w1771 = w679 ~| w1437;
assign w1772 = w681 | w1438;
assign w1773 = w690 | w1438;
assign w1774 = w1030 ~^ w1442;
assign w1775 = w1038 | w1444;
assign w1776 = w1064 ~^ w1445;
assign w1777 = w1034 ~^ w1446;
assign w1778 = w1034 | w1448;
assign w1779 = w1035 ~^ w1449;
assign w1780 = w1035 | w1450;
assign w1781 = w1045 ~^ w1452;
assign w1782 = w1045 | w1453;
assign w1783 = w1069 ~^ w1455;
assign w1784 = w1072 ~^ w1456;
assign w1785 = w1042 | w1457;
assign w1786 = w1076 ~^ w1459;
assign w1787 = w1078 ~^ w1460;
assign w1788 = w354 ~^ w1461;
assign w1789 = w703 | w1462;
assign w1790 = w1036 | w1465;
assign w1791 = w1051 | w1467;
assign w1792 = w1039 ~^ w1474;
assign w1793 = w1039 | w1476;
assign w1794 = w1059 | w1477;
assign w1795 = w358 ~^ w1479;
assign w1796 = w358 | w1480;
assign w1797 = w1055 | w1483;
assign w1798 = w1057 ~^ w1484;
assign w1799 = w1044 | w1485;
assign w1800 = w584 ~| w1487;
assign w1801 = w606 | w1488;
assign w1802 = w605 | w1488;
assign w1803 = w582 ~| w1489;
assign w1804 = w605 | w1489;
assign w1805 = w602 | w1490;
assign w1806 = w591 | w1490;
assign w1807 = w586 ~| w1491;
assign w1808 = w588 | w1492;
assign w1809 = w597 | w1492;
assign w1810 = w967 ~^ w1496;
assign w1811 = w1087 | w1498;
assign w1812 = w1113 ~^ w1499;
assign w1813 = w1083 ~^ w1500;
assign w1814 = w1083 | w1502;
assign w1815 = w1084 ~^ w1503;
assign w1816 = w1084 | w1504;
assign w1817 = w1094 ~^ w1506;
assign w1818 = w1094 | w1507;
assign w1819 = w1118 ~^ w1509;
assign w1820 = w1121 ~^ w1510;
assign w1821 = w1091 | w1511;
assign w1822 = w1125 ~^ w1513;
assign w1823 = w1127 ~^ w1514;
assign w1824 = w378 ~^ w1515;
assign w1825 = w736 | w1516;
assign w1826 = w1085 | w1519;
assign w1827 = w1100 | w1521;
assign w1828 = w1088 ~^ w1528;
assign w1829 = w1088 | w1530;
assign w1830 = w1108 | w1531;
assign w1831 = w382 ~^ w1533;
assign w1832 = w382 | w1534;
assign w1833 = w1104 | w1537;
assign w1834 = w1106 ~^ w1538;
assign w1835 = w1093 | w1539;
assign w1836 = ~w1541;
assign w1837 = w146 & w1546;
assign w1838 = ~w1549;
assign w1839 = ~w1557;
assign w1840 = w181 & w1562;
assign w1841 = ~w1565;
assign w1842 = w168 ~| w1573;
assign w1843 = w822 | w1574;
assign w1844 = w810 | w1574;
assign w1845 = w779 ~| w1575;
assign w1846 = w801 | w1576;
assign w1847 = w800 | w1576;
assign w1848 = w777 ~| w1577;
assign w1849 = w800 | w1577;
assign w1850 = w797 | w1578;
assign w1851 = w786 | w1578;
assign w1852 = w781 ~| w1579;
assign w1853 = w783 | w1580;
assign w1854 = w792 | w1580;
assign w1855 = w1147 ~^ w1584;
assign w1856 = w1155 | w1586;
assign w1857 = w1181 ~^ w1587;
assign w1858 = w1151 ~^ w1588;
assign w1859 = w1151 | w1590;
assign w1860 = w1152 ~^ w1591;
assign w1861 = w1152 | w1592;
assign w1862 = w1162 ~^ w1594;
assign w1863 = w1162 | w1595;
assign w1864 = w1186 ~^ w1597;
assign w1865 = w1189 ~^ w1598;
assign w1866 = w1159 | w1599;
assign w1867 = w1193 ~^ w1601;
assign w1868 = w1195 ~^ w1602;
assign w1869 = w424 ~^ w1603;
assign w1870 = w805 | w1604;
assign w1871 = w1153 | w1607;
assign w1872 = w1168 | w1609;
assign w1873 = w1156 ~^ w1616;
assign w1874 = w1156 | w1618;
assign w1875 = w1176 | w1619;
assign w1876 = w428 ~^ w1621;
assign w1877 = w428 | w1622;
assign w1878 = w1172 | w1625;
assign w1879 = w1174 ~^ w1626;
assign w1880 = w1161 | w1627;
assign w1881 = ~w1629;
assign w1882 = ~w1631;
assign w1883 = w1204 & w1632;
assign w1884 = w864 ~^ w1633;
assign w1885 = w864 | w1633;
assign w1886 = w864 & w1633;
assign w1887 = w846 ^ w1634;
assign w1888 = w846 ~| w1634;
assign w1889 = ~w1637;
assign w1890 = w1636 ~^ w1639;
assign w1891 = w858 & w1639;
assign w1892 = w858 | w1639;
assign w1893 = w1637 ~^ w1640;
assign w1894 = ~w1640;
assign w1895 = ~w1641;
assign w1896 = w13 ^ w1641;
assign w1897 = w1204 & w1642;
assign w1898 = ~w1643;
assign w1899 = w12 ^ w1643;
assign w1900 = ~w1644;
assign w1901 = w14 ^ w1644;
assign w1902 = ~w1645;
assign w1903 = w1225 & w1646;
assign w1904 = w1229 & w1649;
assign w1905 = ~w1650;
assign w1906 = w1233 & w1651;
assign w1907 = w1236 & w1653;
assign w1908 = w1240 & w1656;
assign w1909 = ~w1659;
assign w1910 = w1245 & w1660;
assign w1911 = w1246 & w1661;
assign w1912 = w1248 & w1662;
assign w1913 = ~w1663;
assign w1914 = w1257 & w1664;
assign w1915 = w1260 & w1665;
assign w1916 = ~w1666;
assign w1917 = w1263 & w1667;
assign w1918 = w1264 & w1668;
assign w1919 = w1654 ~^ w1669;
assign w1920 = w1654 ~| w1669;
assign w1921 = w1654 & w1669;
assign w1922 = w1268 & w1670;
assign w1923 = ~w1671;
assign w1924 = ~w1673;
assign w1925 = w1276 & w1674;
assign w1926 = w924 ~^ w1675;
assign w1927 = w924 | w1675;
assign w1928 = w924 & w1675;
assign w1929 = w906 ^ w1676;
assign w1930 = w906 ~| w1676;
assign w1931 = ~w1679;
assign w1932 = w1678 ~^ w1681;
assign w1933 = w918 & w1681;
assign w1934 = w918 | w1681;
assign w1935 = w1679 ~^ w1682;
assign w1936 = ~w1682;
assign w1937 = ~w1683;
assign w1938 = w43 ^ w1683;
assign w1939 = w1276 & w1684;
assign w1940 = ~w1685;
assign w1941 = w42 ^ w1685;
assign w1942 = ~w1686;
assign w1943 = w44 ^ w1686;
assign w1944 = ~w1687;
assign w1945 = w1297 & w1688;
assign w1946 = w1301 & w1691;
assign w1947 = ~w1692;
assign w1948 = w1305 & w1693;
assign w1949 = w1308 & w1695;
assign w1950 = w1312 & w1698;
assign w1951 = ~w1701;
assign w1952 = w1317 & w1702;
assign w1953 = w1318 & w1703;
assign w1954 = w1320 & w1704;
assign w1955 = ~w1705;
assign w1956 = w1329 & w1706;
assign w1957 = w1332 & w1707;
assign w1958 = ~w1708;
assign w1959 = w1335 & w1709;
assign w1960 = w1336 & w1710;
assign w1961 = w1696 ~^ w1711;
assign w1962 = w1696 ~| w1711;
assign w1963 = w1696 & w1711;
assign w1964 = w1340 & w1712;
assign w1965 = ~w1713;
assign w1966 = w1672 ~^ w1714;
assign w1967 = ~w1715;
assign w1968 = w1548 & w1716;
assign w1969 = w1096 ~^ w1717;
assign w1970 = w1096 | w1717;
assign w1971 = w1096 & w1717;
assign w1972 = w966 ^ w1718;
assign w1973 = w966 ~| w1718;
assign w1974 = w1348 & w1719;
assign w1975 = w987 ~^ w1720;
assign w1976 = w987 | w1720;
assign w1977 = w987 & w1720;
assign w1978 = w969 ^ w1721;
assign w1979 = w969 ~| w1721;
assign w1980 = ~w1724;
assign w1981 = w1723 ~^ w1726;
assign w1982 = w981 & w1726;
assign w1983 = w981 | w1726;
assign w1984 = w1724 ~^ w1727;
assign w1985 = ~w1727;
assign w1986 = ~w1728;
assign w1987 = w82 ^ w1728;
assign w1988 = w1348 & w1729;
assign w1989 = ~w1730;
assign w1990 = w81 ^ w1730;
assign w1991 = ~w1731;
assign w1992 = w83 ^ w1731;
assign w1993 = ~w1732;
assign w1994 = w1371 & w1733;
assign w1995 = w1375 & w1736;
assign w1996 = ~w1737;
assign w1997 = w1379 & w1738;
assign w1998 = w1382 & w1740;
assign w1999 = w1386 & w1743;
assign w2000 = ~w1746;
assign w2001 = w1391 & w1747;
assign w2002 = w1392 & w1748;
assign w2003 = w1394 & w1749;
assign w2004 = ~w1750;
assign w2005 = w1403 & w1751;
assign w2006 = w1406 & w1752;
assign w2007 = ~w1753;
assign w2008 = w1409 & w1754;
assign w2009 = w1410 & w1755;
assign w2010 = w1741 ~^ w1756;
assign w2011 = w1741 ~| w1756;
assign w2012 = w1741 & w1756;
assign w2013 = w1414 & w1757;
assign w2014 = ~w1758;
assign w2015 = ~w1759;
assign w2016 = ~w1760;
assign w2017 = w1422 & w1761;
assign w2018 = w1047 ~^ w1762;
assign w2019 = w1047 | w1762;
assign w2020 = w1047 & w1762;
assign w2021 = w1029 ^ w1763;
assign w2022 = w1029 ~| w1763;
assign w2023 = ~w1766;
assign w2024 = w1765 ~^ w1768;
assign w2025 = w1041 & w1768;
assign w2026 = w1041 | w1768;
assign w2027 = w1766 ~^ w1769;
assign w2028 = ~w1769;
assign w2029 = ~w1770;
assign w2030 = w112 ^ w1770;
assign w2031 = w1422 & w1771;
assign w2032 = ~w1772;
assign w2033 = w111 ^ w1772;
assign w2034 = ~w1773;
assign w2035 = w113 ^ w1773;
assign w2036 = ~w1774;
assign w2037 = w1443 & w1775;
assign w2038 = w1447 & w1778;
assign w2039 = ~w1779;
assign w2040 = w1451 & w1780;
assign w2041 = w1454 & w1782;
assign w2042 = w1458 & w1785;
assign w2043 = ~w1788;
assign w2044 = w1463 & w1789;
assign w2045 = w1464 & w1790;
assign w2046 = w1466 & w1791;
assign w2047 = ~w1792;
assign w2048 = w1475 & w1793;
assign w2049 = w1478 & w1794;
assign w2050 = ~w1795;
assign w2051 = w1481 & w1796;
assign w2052 = w1482 & w1797;
assign w2053 = w1783 ~^ w1798;
assign w2054 = w1783 ~| w1798;
assign w2055 = w1783 & w1798;
assign w2056 = w1486 & w1799;
assign w2057 = ~w1802;
assign w2058 = w1801 ~^ w1804;
assign w2059 = w1090 & w1804;
assign w2060 = w1090 | w1804;
assign w2061 = w1802 ~^ w1805;
assign w2062 = ~w1805;
assign w2063 = ~w1806;
assign w2064 = w131 ^ w1806;
assign w2065 = w1548 & w1807;
assign w2066 = ~w1808;
assign w2067 = w130 ^ w1808;
assign w2068 = ~w1809;
assign w2069 = w132 ^ w1809;
assign w2070 = ~w1810;
assign w2071 = w1497 & w1811;
assign w2072 = w1501 & w1814;
assign w2073 = ~w1815;
assign w2074 = w1505 & w1816;
assign w2075 = w1508 & w1818;
assign w2076 = w1512 & w1821;
assign w2077 = ~w1824;
assign w2078 = w1517 & w1825;
assign w2079 = w1518 & w1826;
assign w2080 = w1520 & w1827;
assign w2081 = ~w1828;
assign w2082 = w1529 & w1829;
assign w2083 = w1532 & w1830;
assign w2084 = ~w1831;
assign w2085 = w1535 & w1832;
assign w2086 = w1536 & w1833;
assign w2087 = w1819 ~^ w1834;
assign w2088 = w1819 ~| w1834;
assign w2089 = w1819 & w1834;
assign w2090 = w1540 & w1835;
assign w2091 = ~w1836;
assign w2092 = w1759 ~^ w1837;
assign w2093 = ~w1837;
assign w2094 = ~w1838;
assign w2095 = ~w1839;
assign w2096 = w1672 & w1840;
assign w2097 = w1672 | w1840;
assign w2098 = ~w1841;
assign w2099 = w1564 & w1842;
assign w2100 = w1164 ~^ w1843;
assign w2101 = w1164 | w1843;
assign w2102 = w1164 & w1843;
assign w2103 = w1146 ^ w1844;
assign w2104 = w1146 ~| w1844;
assign w2105 = ~w1847;
assign w2106 = w1846 ~^ w1849;
assign w2107 = w1158 & w1849;
assign w2108 = w1158 | w1849;
assign w2109 = w1847 ~^ w1850;
assign w2110 = ~w1850;
assign w2111 = ~w1851;
assign w2112 = w166 ^ w1851;
assign w2113 = w1564 & w1852;
assign w2114 = ~w1853;
assign w2115 = w165 ^ w1853;
assign w2116 = ~w1854;
assign w2117 = w167 ^ w1854;
assign w2118 = ~w1855;
assign w2119 = w1585 & w1856;
assign w2120 = w1589 & w1859;
assign w2121 = ~w1860;
assign w2122 = w1593 & w1861;
assign w2123 = w1596 & w1863;
assign w2124 = w1600 & w1866;
assign w2125 = ~w1869;
assign w2126 = w1605 & w1870;
assign w2127 = w1606 & w1871;
assign w2128 = w1608 & w1872;
assign w2129 = ~w1873;
assign w2130 = w1617 & w1874;
assign w2131 = w1620 & w1875;
assign w2132 = ~w1876;
assign w2133 = w1623 & w1877;
assign w2134 = w1624 & w1878;
assign w2135 = w1864 ~^ w1879;
assign w2136 = w1864 ~| w1879;
assign w2137 = w1864 & w1879;
assign w2138 = w1628 & w1880;
assign w2139 = w1635 & w1881;
assign w2140 = w1638 & w1882;
assign w2141 = in5[0] ~^ w1883;
assign w2142 = w1883 & in5[0];
assign w2143 = w854 ~^ w1884;
assign w2144 = w854 | w1886;
assign w2145 = w1212 & w1887;
assign w2146 = w1203 & w1888;
assign w2147 = w858 ~^ w1890;
assign w2148 = w1636 | w1891;
assign w2149 = ~w1893;
assign w2150 = w1889 & w1894;
assign w2151 = w13 & w1895;
assign w2152 = w12 & w1898;
assign w2153 = w1221 ^ w1899;
assign w2154 = w1222 ~| w1899;
assign w2155 = w14 & w1900;
assign w2156 = w1647 ~^ w1903;
assign w2157 = w1901 ~^ w1906;
assign w2158 = w1901 | w1906;
assign w2159 = w1901 & w1906;
assign w2160 = w207 ~^ w1907;
assign w2161 = w483 | w1907;
assign w2162 = ~w1907;
assign w2163 = w888 ~^ w1908;
assign w2164 = w888 & w1908;
assign w2165 = w888 | w1908;
assign w2166 = w1657 ~^ w1912;
assign w2167 = w1657 ~| w1912;
assign w2168 = w1657 & w1912;
assign w2169 = w1253 ^ w1915;
assign w2170 = w1254 ~| w1915;
assign w2171 = w1645 ~^ w1917;
assign w2172 = w1645 ~| w1917;
assign w2173 = ~w1917;
assign w2174 = w1250 ~^ w1918;
assign w2175 = w1252 | w1918;
assign w2176 = w1910 ~^ w1919;
assign w2177 = w1910 ~| w1921;
assign w2178 = w1911 ~^ w1922;
assign w2179 = w1911 & w1922;
assign w2180 = w1911 | w1922;
assign w2181 = w1677 & w1923;
assign w2182 = w1680 & w1924;
assign w2183 = ~w1925;
assign w2184 = w914 ~^ w1926;
assign w2185 = w914 | w1928;
assign w2186 = w1284 & w1929;
assign w2187 = w1275 & w1930;
assign w2188 = w918 ~^ w1932;
assign w2189 = w1678 | w1933;
assign w2190 = ~w1935;
assign w2191 = w1931 & w1936;
assign w2192 = w43 & w1937;
assign w2193 = w42 & w1940;
assign w2194 = w1293 ^ w1941;
assign w2195 = w1294 ~| w1941;
assign w2196 = w44 & w1942;
assign w2197 = w1689 ~^ w1945;
assign w2198 = w1943 ~^ w1948;
assign w2199 = w1943 | w1948;
assign w2200 = w1943 & w1948;
assign w2201 = w251 ~^ w1949;
assign w2202 = w548 | w1949;
assign w2203 = ~w1949;
assign w2204 = w948 ~^ w1950;
assign w2205 = w948 & w1950;
assign w2206 = w948 | w1950;
assign w2207 = w1699 ~^ w1954;
assign w2208 = w1699 ~| w1954;
assign w2209 = w1699 & w1954;
assign w2210 = w1325 ^ w1957;
assign w2211 = w1326 ~| w1957;
assign w2212 = w1687 ~^ w1959;
assign w2213 = w1687 ~| w1959;
assign w2214 = ~w1959;
assign w2215 = w1322 ~^ w1960;
assign w2216 = w1324 | w1960;
assign w2217 = w1952 ~^ w1961;
assign w2218 = w1952 ~| w1963;
assign w2219 = w1953 ~^ w1964;
assign w2220 = w1953 & w1964;
assign w2221 = w1953 | w1964;
assign w2222 = w1722 & w1965;
assign w2223 = w1840 ~^ w1966;
assign w2224 = w1725 & w1967;
assign w2225 = ~w1968;
assign w2226 = w1086 ~^ w1969;
assign w2227 = w1086 | w1971;
assign w2228 = w1556 & w1972;
assign w2229 = w1547 & w1973;
assign w2230 = w1925 ~| w1974;
assign w2231 = ~w1974;
assign w2232 = w977 ~^ w1975;
assign w2233 = w977 | w1977;
assign w2234 = w1356 & w1978;
assign w2235 = w1347 & w1979;
assign w2236 = w981 ~^ w1981;
assign w2237 = w1723 | w1982;
assign w2238 = ~w1984;
assign w2239 = w1980 & w1985;
assign w2240 = w82 & w1986;
assign w2241 = w81 & w1989;
assign w2242 = w1367 ^ w1990;
assign w2243 = w1368 ~| w1990;
assign w2244 = w83 & w1991;
assign w2245 = w1734 ~^ w1994;
assign w2246 = w1992 ~^ w1997;
assign w2247 = w1992 | w1997;
assign w2248 = w1992 & w1997;
assign w2249 = w313 ~^ w1998;
assign w2250 = w641 | w1998;
assign w2251 = ~w1998;
assign w2252 = w1011 ~^ w1999;
assign w2253 = w1011 & w1999;
assign w2254 = w1011 | w1999;
assign w2255 = w1744 ~^ w2003;
assign w2256 = w1744 ~| w2003;
assign w2257 = w1744 & w2003;
assign w2258 = w1399 ^ w2006;
assign w2259 = w1400 ~| w2006;
assign w2260 = w1732 ~^ w2008;
assign w2261 = w1732 ~| w2008;
assign w2262 = ~w2008;
assign w2263 = w1396 ~^ w2009;
assign w2264 = w1398 | w2009;
assign w2265 = w2001 ~^ w2010;
assign w2266 = w2001 ~| w2012;
assign w2267 = w2002 ~^ w2013;
assign w2268 = w2002 & w2013;
assign w2269 = w2002 | w2013;
assign w2270 = w1764 & w2014;
assign w2271 = w1767 & w2016;
assign w2272 = w1968 & w2017;
assign w2273 = w1037 ~^ w2018;
assign w2274 = w1037 | w2020;
assign w2275 = w1430 & w2021;
assign w2276 = w1421 & w2022;
assign w2277 = w1041 ~^ w2024;
assign w2278 = w1765 | w2025;
assign w2279 = ~w2027;
assign w2280 = w2023 & w2028;
assign w2281 = w112 & w2029;
assign w2282 = w2031 ~^ in5[2];
assign w2283 = ~w2031;
assign w2284 = w111 & w2032;
assign w2285 = w1439 ^ w2033;
assign w2286 = w1440 ~| w2033;
assign w2287 = w113 & w2034;
assign w2288 = w1776 ~^ w2037;
assign w2289 = w2035 ~^ w2040;
assign w2290 = w2035 | w2040;
assign w2291 = w2035 & w2040;
assign w2292 = w357 ~^ w2041;
assign w2293 = w706 | w2041;
assign w2294 = ~w2041;
assign w2295 = w1071 ~^ w2042;
assign w2296 = w1071 & w2042;
assign w2297 = w1071 | w2042;
assign w2298 = w1786 ~^ w2046;
assign w2299 = w1786 ~| w2046;
assign w2300 = w1786 & w2046;
assign w2301 = w1471 ^ w2049;
assign w2302 = w1472 ~| w2049;
assign w2303 = w1774 ~^ w2051;
assign w2304 = w1774 ~| w2051;
assign w2305 = ~w2051;
assign w2306 = w1468 ~^ w2052;
assign w2307 = w1470 | w2052;
assign w2308 = w2044 ~^ w2053;
assign w2309 = w2044 ~| w2055;
assign w2310 = w2045 ~^ w2056;
assign w2311 = w2045 & w2056;
assign w2312 = w2045 | w2056;
assign w2313 = w1090 ~^ w2058;
assign w2314 = w1801 | w2059;
assign w2315 = ~w2061;
assign w2316 = w2057 & w2062;
assign w2317 = w131 & w2063;
assign w2318 = w130 & w2066;
assign w2319 = w1493 ^ w2067;
assign w2320 = w1494 ~| w2067;
assign w2321 = w132 & w2068;
assign w2322 = w1812 ~^ w2071;
assign w2323 = w2069 ~^ w2074;
assign w2324 = w2069 | w2074;
assign w2325 = w2069 & w2074;
assign w2326 = w381 ~^ w2075;
assign w2327 = w739 | w2075;
assign w2328 = ~w2075;
assign w2329 = w1120 ~^ w2076;
assign w2330 = w1120 & w2076;
assign w2331 = w1120 | w2076;
assign w2332 = w1822 ~^ w2080;
assign w2333 = w1822 ~| w2080;
assign w2334 = w1822 & w2080;
assign w2335 = w1525 ^ w2083;
assign w2336 = w1526 ~| w2083;
assign w2337 = w1810 ~^ w2085;
assign w2338 = w1810 ~| w2085;
assign w2339 = ~w2085;
assign w2340 = w1522 ~^ w2086;
assign w2341 = w1524 | w2086;
assign w2342 = w2078 ~^ w2087;
assign w2343 = w2078 ~| w2089;
assign w2344 = w2079 ~^ w2090;
assign w2345 = w2079 & w2090;
assign w2346 = w2079 | w2090;
assign w2347 = w1800 & w2091;
assign w2348 = w1630 ~^ w2092;
assign w2349 = w2015 | w2093;
assign w2350 = w1803 & w2094;
assign w2351 = w1845 & w2095;
assign w2352 = w1714 & w2097;
assign w2353 = w1848 & w2098;
assign w2354 = w1974 ~^ w2099;
assign w2355 = ~w2099;
assign w2356 = w1154 ~^ w2100;
assign w2357 = w1154 | w2102;
assign w2358 = w1572 & w2103;
assign w2359 = w1563 & w2104;
assign w2360 = w1158 ~^ w2106;
assign w2361 = w1846 | w2107;
assign w2362 = ~w2109;
assign w2363 = w2105 & w2110;
assign w2364 = w166 & w2111;
assign w2365 = w165 & w2114;
assign w2366 = w1581 ^ w2115;
assign w2367 = w1582 ~| w2115;
assign w2368 = w167 & w2116;
assign w2369 = w1857 ~^ w2119;
assign w2370 = w2117 ~^ w2122;
assign w2371 = w2117 | w2122;
assign w2372 = w2117 & w2122;
assign w2373 = w427 ~^ w2123;
assign w2374 = w808 | w2123;
assign w2375 = ~w2123;
assign w2376 = w1188 ~^ w2124;
assign w2377 = w1188 & w2124;
assign w2378 = w1188 | w2124;
assign w2379 = w1867 ~^ w2128;
assign w2380 = w1867 ~| w2128;
assign w2381 = w1867 & w2128;
assign w2382 = w1613 ^ w2131;
assign w2383 = w1614 ~| w2131;
assign w2384 = w1855 ~^ w2133;
assign w2385 = w1855 ~| w2133;
assign w2386 = ~w2133;
assign w2387 = w1610 ~^ w2134;
assign w2388 = w1612 | w2134;
assign w2389 = w2126 ~^ w2135;
assign w2390 = w2126 ~| w2137;
assign w2391 = w2127 ~^ w2138;
assign w2392 = w2127 & w2138;
assign w2393 = w2127 | w2138;
assign w2394 = in5[1] ~| w2139;
assign w2395 = ~w2139;
assign w2396 = ~w2141;
assign w2397 = ~w2142;
assign w2398 = w1885 & w2144;
assign w2399 = w1939 ~^ w2145;
assign w2400 = w1939 & w2145;
assign w2401 = w1939 ~| w2145;
assign w2402 = w1892 & w2148;
assign w2403 = w502 ~^ w2150;
assign w2404 = w221 & w2150;
assign w2405 = w498 ~^ w2151;
assign w2406 = w24 ~| w2151;
assign w2407 = ~w2151;
assign w2408 = w1896 ~^ w2152;
assign w2409 = ~w2152;
assign w2410 = w1211 & w2153;
assign w2411 = w1223 | w2154;
assign w2412 = w1893 ~^ w2155;
assign w2413 = w2149 ~| w2155;
assign w2414 = ~w2155;
assign w2415 = w1648 ~^ w2157;
assign w2416 = w1648 | w2159;
assign w2417 = w1658 ~^ w2160;
assign w2418 = w207 ~| w2162;
assign w2419 = w1655 ~^ w2163;
assign w2420 = w1655 | w2164;
assign w2421 = w1199 & w2169;
assign w2422 = w1255 | w2170;
assign w2423 = w1902 | w2173;
assign w2424 = w2156 ~^ w2174;
assign w2425 = w1647 | w2174;
assign w2426 = w1647 & w2174;
assign w2427 = w1251 & w2175;
assign w2428 = w1920 | w2177;
assign w2429 = w2147 ~^ w2178;
assign w2430 = w2147 | w2179;
assign w2431 = w1927 & w2185;
assign w2432 = w1934 & w2189;
assign w2433 = w567 ~^ w2191;
assign w2434 = w265 & w2191;
assign w2435 = w563 ~^ w2192;
assign w2436 = w54 ~| w2192;
assign w2437 = ~w2192;
assign w2438 = w1938 ~^ w2193;
assign w2439 = ~w2193;
assign w2440 = w1283 & w2194;
assign w2441 = w1295 | w2195;
assign w2442 = w1935 ~^ w2196;
assign w2443 = w2190 ~| w2196;
assign w2444 = ~w2196;
assign w2445 = w1690 ~^ w2198;
assign w2446 = w1690 | w2200;
assign w2447 = w1700 ~^ w2201;
assign w2448 = w251 ~| w2203;
assign w2449 = w1697 ~^ w2204;
assign w2450 = w1697 | w2205;
assign w2451 = w1271 & w2210;
assign w2452 = w1327 | w2211;
assign w2453 = w1944 | w2214;
assign w2454 = w2197 ~^ w2215;
assign w2455 = w1689 | w2215;
assign w2456 = w1689 & w2215;
assign w2457 = w1323 & w2216;
assign w2458 = w1962 | w2218;
assign w2459 = w2188 ~^ w2219;
assign w2460 = w2188 | w2220;
assign w2461 = w2181 ~^ w2222;
assign w2462 = w2181 & w2222;
assign w2463 = w2181 | w2222;
assign w2464 = w2017 ~^ w2225;
assign w2465 = w1970 & w2227;
assign w2466 = w2113 ~^ w2228;
assign w2467 = w2113 | w2228;
assign w2468 = w2113 & w2228;
assign w2469 = w2183 | w2231;
assign w2470 = w1976 & w2233;
assign w2471 = w1897 ~^ w2234;
assign w2472 = w1897 | w2234;
assign w2473 = w1897 & w2234;
assign w2474 = w2229 ~^ w2235;
assign w2475 = w2229 | w2235;
assign w2476 = w2229 & w2235;
assign w2477 = w1983 & w2237;
assign w2478 = w660 ~^ w2239;
assign w2479 = w327 & w2239;
assign w2480 = w656 ~^ w2240;
assign w2481 = w93 ~| w2240;
assign w2482 = ~w2240;
assign w2483 = w1987 ~^ w2241;
assign w2484 = ~w2241;
assign w2485 = w1355 & w2242;
assign w2486 = w1369 | w2243;
assign w2487 = w1984 ~^ w2244;
assign w2488 = w2238 ~| w2244;
assign w2489 = ~w2244;
assign w2490 = w1735 ~^ w2246;
assign w2491 = w1735 | w2248;
assign w2492 = w1745 ~^ w2249;
assign w2493 = w313 ~| w2251;
assign w2494 = w1742 ~^ w2252;
assign w2495 = w1742 | w2253;
assign w2496 = w1343 & w2258;
assign w2497 = w1401 | w2259;
assign w2498 = w1993 | w2262;
assign w2499 = w2245 ~^ w2263;
assign w2500 = w1734 | w2263;
assign w2501 = w1734 & w2263;
assign w2502 = w1397 & w2264;
assign w2503 = w2011 | w2266;
assign w2504 = w2236 ~^ w2267;
assign w2505 = w2236 | w2268;
assign w2506 = w2270 ~^ in5[1];
assign w2507 = ~w2270;
assign w2508 = w2142 ~^ w2271;
assign w2509 = w2019 & w2274;
assign w2510 = w2186 ~^ w2275;
assign w2511 = w2186 & w2275;
assign w2512 = w2186 | w2275;
assign w2513 = w2276 ~^ in5[3];
assign w2514 = ~w2276;
assign w2515 = w2026 & w2278;
assign w2516 = w725 ~^ w2280;
assign w2517 = w371 & w2280;
assign w2518 = w721 ~^ w2281;
assign w2519 = w123 ~| w2281;
assign w2520 = ~w2281;
assign w2521 = w151 | w2283;
assign w2522 = w2030 ~^ w2284;
assign w2523 = ~w2284;
assign w2524 = w1429 & w2285;
assign w2525 = w1441 | w2286;
assign w2526 = w2027 ~^ w2287;
assign w2527 = w2279 ~| w2287;
assign w2528 = ~w2287;
assign w2529 = w1777 ~^ w2289;
assign w2530 = w1777 | w2291;
assign w2531 = w1787 ~^ w2292;
assign w2532 = w357 ~| w2294;
assign w2533 = w1784 ~^ w2295;
assign w2534 = w1784 | w2296;
assign w2535 = w1417 & w2301;
assign w2536 = w1473 | w2302;
assign w2537 = w2036 | w2305;
assign w2538 = w2288 ~^ w2306;
assign w2539 = w1776 | w2306;
assign w2540 = w1776 & w2306;
assign w2541 = w1469 & w2307;
assign w2542 = w2054 | w2309;
assign w2543 = w2277 ~^ w2310;
assign w2544 = w2277 | w2311;
assign w2545 = w2060 & w2314;
assign w2546 = w758 ~^ w2316;
assign w2547 = w395 & w2316;
assign w2548 = w754 ~^ w2317;
assign w2549 = w142 ~| w2317;
assign w2550 = ~w2317;
assign w2551 = w2064 ~^ w2318;
assign w2552 = ~w2318;
assign w2553 = w1555 & w2319;
assign w2554 = w1495 | w2320;
assign w2555 = w2061 ~^ w2321;
assign w2556 = w2315 ~| w2321;
assign w2557 = ~w2321;
assign w2558 = w1813 ~^ w2323;
assign w2559 = w1813 | w2325;
assign w2560 = w1823 ~^ w2326;
assign w2561 = w381 ~| w2328;
assign w2562 = w1820 ~^ w2329;
assign w2563 = w1820 | w2330;
assign w2564 = w1543 & w2335;
assign w2565 = w1527 | w2336;
assign w2566 = w2070 | w2339;
assign w2567 = w2322 ~^ w2340;
assign w2568 = w1812 | w2340;
assign w2569 = w1812 & w2340;
assign w2570 = w1523 & w2341;
assign w2571 = w2088 | w2343;
assign w2572 = w2313 ~^ w2344;
assign w2573 = w2313 | w2345;
assign w2574 = ~w2349;
assign w2575 = w2347 ~^ w2351;
assign w2576 = w2347 | w2351;
assign w2577 = w2347 & w2351;
assign w2578 = w2096 | w2352;
assign w2579 = w2224 ~^ w2353;
assign w2580 = w2140 & w2353;
assign w2581 = w2140 | w2353;
assign w2582 = w1925 ~^ w2354;
assign w2583 = w2230 | w2355;
assign w2584 = w2101 & w2357;
assign w2585 = w2146 ~^ w2359;
assign w2586 = w2146 & w2359;
assign w2587 = w2146 | w2359;
assign w2588 = w2108 & w2361;
assign w2589 = w827 ~^ w2363;
assign w2590 = w441 & w2363;
assign w2591 = w823 ~^ w2364;
assign w2592 = w177 ~| w2364;
assign w2593 = ~w2364;
assign w2594 = w2112 ~^ w2365;
assign w2595 = ~w2365;
assign w2596 = w1571 & w2366;
assign w2597 = w1583 | w2367;
assign w2598 = w2109 ~^ w2368;
assign w2599 = w2362 ~| w2368;
assign w2600 = ~w2368;
assign w2601 = w1858 ~^ w2370;
assign w2602 = w1858 | w2372;
assign w2603 = w1868 ~^ w2373;
assign w2604 = w427 ~| w2375;
assign w2605 = w1865 ~^ w2376;
assign w2606 = w1865 | w2377;
assign w2607 = w1559 & w2382;
assign w2608 = w1615 | w2383;
assign w2609 = w2118 | w2386;
assign w2610 = w2369 ~^ w2387;
assign w2611 = w1857 | w2387;
assign w2612 = w1857 & w2387;
assign w2613 = w1611 & w2388;
assign w2614 = w2136 | w2390;
assign w2615 = w2360 ~^ w2391;
assign w2616 = w2360 | w2392;
assign w2617 = w150 | w2395;
assign w2618 = w1650 ~^ w2398;
assign w2619 = w1650 ~| w2398;
assign w2620 = ~w2398;
assign w2621 = w2282 ~^ w2399;
assign w2622 = w2282 ~| w2401;
assign w2623 = w1914 ~^ w2402;
assign w2624 = w1914 | w2402;
assign w2625 = w1914 & w2402;
assign w2626 = w1663 ~^ w2403;
assign w2627 = w1913 ~| w2403;
assign w2628 = ~w2403;
assign w2629 = w503 | w2404;
assign w2630 = w205 | w2406;
assign w2631 = w218 | w2407;
assign w2632 = w2143 ~^ w2408;
assign w2633 = w1896 & w2409;
assign w2634 = w1896 ~| w2409;
assign w2635 = ~w2410;
assign w2636 = w1199 & w2411;
assign w2637 = w1904 ~^ w2412;
assign w2638 = w1904 | w2413;
assign w2639 = w1893 | w2414;
assign w2640 = w2158 & w2416;
assign w2641 = w2171 ~^ w2417;
assign w2642 = w1658 | w2418;
assign w2643 = w2165 & w2420;
assign w2644 = w1210 & w2422;
assign w2645 = w2417 & w2423;
assign w2646 = ~w2424;
assign w2647 = w1903 | w2426;
assign w2648 = w2419 ~^ w2427;
assign w2649 = w2419 ~| w2427;
assign w2650 = w2419 & w2427;
assign w2651 = ~w2428;
assign w2652 = ~w2429;
assign w2653 = w2180 & w2430;
assign w2654 = w1692 ~^ w2431;
assign w2655 = w1692 ~| w2431;
assign w2656 = ~w2431;
assign w2657 = w1956 ~^ w2432;
assign w2658 = w1956 | w2432;
assign w2659 = w1956 & w2432;
assign w2660 = w1705 ~^ w2433;
assign w2661 = w1955 ~| w2433;
assign w2662 = ~w2433;
assign w2663 = w568 | w2434;
assign w2664 = w249 | w2436;
assign w2665 = w262 | w2437;
assign w2666 = w2184 ~^ w2438;
assign w2667 = w1938 & w2439;
assign w2668 = w1938 ~| w2439;
assign w2669 = w1271 & w2441;
assign w2670 = w1946 ~^ w2442;
assign w2671 = w1946 | w2443;
assign w2672 = w1935 | w2444;
assign w2673 = w2199 & w2446;
assign w2674 = w2212 ~^ w2447;
assign w2675 = w1700 | w2448;
assign w2676 = w2206 & w2450;
assign w2677 = w1282 & w2452;
assign w2678 = w2447 & w2453;
assign w2679 = ~w2454;
assign w2680 = w1945 | w2456;
assign w2681 = w2449 ~^ w2457;
assign w2682 = w2449 ~| w2457;
assign w2683 = w2449 & w2457;
assign w2684 = ~w2458;
assign w2685 = ~w2459;
assign w2686 = w2221 & w2460;
assign w2687 = w2182 ~^ w2461;
assign w2688 = w2182 & w2463;
assign w2689 = w1815 ~^ w2465;
assign w2690 = w1815 ~| w2465;
assign w2691 = ~w2465;
assign w2692 = w1988 ~^ w2466;
assign w2693 = w1988 & w2467;
assign w2694 = w1737 ~^ w2470;
assign w2695 = w1737 ~| w2470;
assign w2696 = ~w2470;
assign w2697 = w2358 ~^ w2471;
assign w2698 = w2358 & w2472;
assign w2699 = w2440 ^ w2474;
assign w2700 = w2440 & w2475;
assign w2701 = w2005 ~^ w2477;
assign w2702 = w2005 | w2477;
assign w2703 = w2005 & w2477;
assign w2704 = w1750 ~^ w2478;
assign w2705 = w2004 ~| w2478;
assign w2706 = ~w2478;
assign w2707 = w661 | w2479;
assign w2708 = w311 | w2481;
assign w2709 = w324 | w2482;
assign w2710 = w2232 ~^ w2483;
assign w2711 = w1987 & w2484;
assign w2712 = w1987 ~| w2484;
assign w2713 = w1343 & w2486;
assign w2714 = w1995 ~^ w2487;
assign w2715 = w1995 | w2488;
assign w2716 = w1984 | w2489;
assign w2717 = w2247 & w2491;
assign w2718 = w2260 ~^ w2492;
assign w2719 = w1745 | w2493;
assign w2720 = w2254 & w2495;
assign w2721 = w2451 ~^ w2496;
assign w2722 = w2451 & w2496;
assign w2723 = w2451 | w2496;
assign w2724 = w1354 & w2497;
assign w2725 = w2492 & w2498;
assign w2726 = ~w2499;
assign w2727 = w1994 | w2501;
assign w2728 = w2494 ~^ w2502;
assign w2729 = w2494 ~| w2502;
assign w2730 = w2494 & w2502;
assign w2731 = ~w2503;
assign w2732 = ~w2504;
assign w2733 = w2269 & w2505;
assign w2734 = w2139 ^ w2506;
assign w2735 = w2394 | w2507;
assign w2736 = w1779 ~^ w2509;
assign w2737 = w1779 ~| w2509;
assign w2738 = ~w2509;
assign w2739 = w2065 ^ w2510;
assign w2740 = w2065 & w2512;
assign w2741 = w152 | w2514;
assign w2742 = w2048 ~^ w2515;
assign w2743 = w2048 | w2515;
assign w2744 = w2048 & w2515;
assign w2745 = w1792 ~^ w2516;
assign w2746 = w2047 ~| w2516;
assign w2747 = ~w2516;
assign w2748 = w726 | w2517;
assign w2749 = w355 | w2519;
assign w2750 = w368 | w2520;
assign w2751 = ~w2521;
assign w2752 = w2273 ~^ w2522;
assign w2753 = w2030 & w2523;
assign w2754 = w2030 ~| w2523;
assign w2755 = w2485 ~^ w2524;
assign w2756 = w2485 & w2524;
assign w2757 = w2485 | w2524;
assign w2758 = w1417 & w2525;
assign w2759 = w2038 ~^ w2526;
assign w2760 = w2038 | w2527;
assign w2761 = w2027 | w2528;
assign w2762 = w2290 & w2530;
assign w2763 = w2303 ~^ w2531;
assign w2764 = w1787 | w2532;
assign w2765 = w2297 & w2534;
assign w2766 = ~w2535;
assign w2767 = w1428 & w2536;
assign w2768 = w2531 & w2537;
assign w2769 = ~w2538;
assign w2770 = w2037 | w2540;
assign w2771 = w2533 ~^ w2541;
assign w2772 = w2533 ~| w2541;
assign w2773 = w2533 & w2541;
assign w2774 = ~w2542;
assign w2775 = ~w2543;
assign w2776 = w2312 & w2544;
assign w2777 = w2082 ~^ w2545;
assign w2778 = w2082 | w2545;
assign w2779 = w2082 & w2545;
assign w2780 = w1828 ~^ w2546;
assign w2781 = w2081 ~| w2546;
assign w2782 = ~w2546;
assign w2783 = w759 | w2547;
assign w2784 = w379 | w2549;
assign w2785 = w392 | w2550;
assign w2786 = w2226 ~^ w2551;
assign w2787 = w2064 & w2552;
assign w2788 = w2064 ~| w2552;
assign w2789 = w1543 & w2554;
assign w2790 = w2072 ~^ w2555;
assign w2791 = w2072 | w2556;
assign w2792 = w2061 | w2557;
assign w2793 = w2324 & w2559;
assign w2794 = w2337 ~^ w2560;
assign w2795 = w1823 | w2561;
assign w2796 = w2331 & w2563;
assign w2797 = w2535 ~^ w2564;
assign w2798 = ~w2564;
assign w2799 = w1554 & w2565;
assign w2800 = w2560 & w2566;
assign w2801 = ~w2567;
assign w2802 = w2071 | w2569;
assign w2803 = w2562 ~^ w2570;
assign w2804 = w2562 ~| w2570;
assign w2805 = w2562 & w2570;
assign w2806 = ~w2571;
assign w2807 = ~w2572;
assign w2808 = w2346 & w2573;
assign w2809 = w2350 ~^ w2575;
assign w2810 = w2350 & w2576;
assign w2811 = w2140 ~^ w2579;
assign w2812 = w2224 & w2581;
assign w2813 = w2396 ~^ w2582;
assign w2814 = w2464 & w2582;
assign w2815 = w2464 | w2582;
assign w2816 = w2469 & w2583;
assign w2817 = w1860 ~^ w2584;
assign w2818 = w1860 ~| w2584;
assign w2819 = ~w2584;
assign w2820 = w2187 ~^ w2585;
assign w2821 = w2187 & w2587;
assign w2822 = w2130 ~^ w2588;
assign w2823 = w2130 | w2588;
assign w2824 = w2130 & w2588;
assign w2825 = w1873 ~^ w2589;
assign w2826 = w2129 ~| w2589;
assign w2827 = ~w2589;
assign w2828 = w828 | w2590;
assign w2829 = w425 | w2592;
assign w2830 = w438 | w2593;
assign w2831 = w2356 ~^ w2594;
assign w2832 = w2112 & w2595;
assign w2833 = w2112 ~| w2595;
assign w2834 = w2410 ~^ w2596;
assign w2835 = w2410 ~| w2596;
assign w2836 = ~w2596;
assign w2837 = w1559 & w2597;
assign w2838 = w2120 ~^ w2598;
assign w2839 = w2120 | w2599;
assign w2840 = w2109 | w2600;
assign w2841 = w2371 & w2602;
assign w2842 = w2384 ~^ w2603;
assign w2843 = w1868 | w2604;
assign w2844 = w2378 & w2606;
assign w2845 = w1570 & w2608;
assign w2846 = w2603 & w2609;
assign w2847 = ~w2610;
assign w2848 = w2119 | w2612;
assign w2849 = w2605 ~^ w2613;
assign w2850 = w2605 ~| w2613;
assign w2851 = w2605 & w2613;
assign w2852 = ~w2614;
assign w2853 = ~w2615;
assign w2854 = w2393 & w2616;
assign w2855 = w2405 ~^ w2618;
assign w2856 = w1905 | w2620;
assign w2857 = w2400 | w2622;
assign w2858 = w1652 ~^ w2623;
assign w2859 = w1652 | w2625;
assign w2860 = w1663 | w2628;
assign w2861 = w1666 ~^ w2629;
assign w2862 = w1916 ~| w2629;
assign w2863 = ~w2629;
assign w2864 = w2630 & w2631;
assign w2865 = w1207 & w2632;
assign w2866 = w2143 ~| w2633;
assign w2867 = in5[4] & w2636;
assign w2868 = in5[4] | w2636;
assign w2869 = ~w2637;
assign w2870 = w2638 & w2639;
assign w2871 = w2637 ~^ w2640;
assign w2872 = ~w2641;
assign w2873 = w2161 & w2642;
assign w2874 = w2166 ^ w2643;
assign w2875 = w2168 ~| w2643;
assign w2876 = w2172 | w2645;
assign w2877 = w2425 & w2647;
assign w2878 = w2429 ~^ w2651;
assign w2879 = w2429 ~| w2651;
assign w2880 = w2428 | w2652;
assign w2881 = w2435 ~^ w2654;
assign w2882 = w1947 | w2656;
assign w2883 = w1694 ~^ w2657;
assign w2884 = w1694 | w2659;
assign w2885 = w1705 | w2662;
assign w2886 = w1708 ~^ w2663;
assign w2887 = w1958 ~| w2663;
assign w2888 = ~w2663;
assign w2889 = w2664 & w2665;
assign w2890 = w1279 & w2666;
assign w2891 = w2184 ~| w2667;
assign w2892 = ~w2669;
assign w2893 = ~w2670;
assign w2894 = w2671 & w2672;
assign w2895 = w2670 ~^ w2673;
assign w2896 = ~w2674;
assign w2897 = w2202 & w2675;
assign w2898 = w2207 ^ w2676;
assign w2899 = w2209 ~| w2676;
assign w2900 = w2348 ~^ w2677;
assign w2901 = w1630 & w2677;
assign w2902 = w1630 ~| w2677;
assign w2903 = w2213 | w2678;
assign w2904 = w2455 & w2680;
assign w2905 = w2459 ~^ w2684;
assign w2906 = w2459 ~| w2684;
assign w2907 = w2458 | w2685;
assign w2908 = w2272 & w2687;
assign w2909 = w2272 ~| w2687;
assign w2910 = w2462 | w2688;
assign w2911 = w2548 ~^ w2689;
assign w2912 = w2073 | w2691;
assign w2913 = w2621 ~^ w2692;
assign w2914 = ~w2692;
assign w2915 = w2468 | w2693;
assign w2916 = w2480 ~^ w2694;
assign w2917 = w1996 | w2696;
assign w2918 = w2473 | w2698;
assign w2919 = w2476 | w2700;
assign w2920 = w1739 ~^ w2701;
assign w2921 = w1739 | w2703;
assign w2922 = w1750 | w2706;
assign w2923 = w1753 ~^ w2707;
assign w2924 = w2007 ~| w2707;
assign w2925 = ~w2707;
assign w2926 = w2708 & w2709;
assign w2927 = w1351 & w2710;
assign w2928 = w2232 ~| w2711;
assign w2929 = ~w2714;
assign w2930 = w2715 & w2716;
assign w2931 = w2714 ~^ w2717;
assign w2932 = ~w2718;
assign w2933 = w2250 & w2719;
assign w2934 = w2255 ^ w2720;
assign w2935 = w2257 ~| w2720;
assign w2936 = w2607 ~^ w2721;
assign w2937 = w2607 & w2723;
assign w2938 = w2644 ~^ w2724;
assign w2939 = w2261 | w2725;
assign w2940 = w2500 & w2727;
assign w2941 = w2504 ~^ w2731;
assign w2942 = w2504 ~| w2731;
assign w2943 = w2503 | w2732;
assign w2944 = w2617 & w2735;
assign w2945 = w2518 ~^ w2736;
assign w2946 = w2039 | w2738;
assign w2947 = w2511 | w2740;
assign w2948 = w2669 ~^ w2741;
assign w2949 = ~w2741;
assign w2950 = w1781 ~^ w2742;
assign w2951 = w1781 | w2744;
assign w2952 = w1792 | w2747;
assign w2953 = w1795 ~^ w2748;
assign w2954 = w2050 ~| w2748;
assign w2955 = ~w2748;
assign w2956 = w2749 & w2750;
assign w2957 = w1425 & w2752;
assign w2958 = w2273 ~| w2753;
assign w2959 = w2553 ~^ w2755;
assign w2960 = w2553 & w2757;
assign w2961 = w2758 ~^ in5[4];
assign w2962 = ~w2759;
assign w2963 = w2760 & w2761;
assign w2964 = w2759 ~^ w2762;
assign w2965 = ~w2763;
assign w2966 = w2293 & w2764;
assign w2967 = w2298 ^ w2765;
assign w2968 = w2300 ~| w2765;
assign w2969 = w2724 | w2767;
assign w2970 = w2724 & w2767;
assign w2971 = w2304 | w2768;
assign w2972 = w2539 & w2770;
assign w2973 = w2543 ~^ w2774;
assign w2974 = w2543 ~| w2774;
assign w2975 = w2542 | w2775;
assign w2976 = w1817 ~^ w2777;
assign w2977 = w1817 | w2779;
assign w2978 = w1828 | w2782;
assign w2979 = w1831 ~^ w2783;
assign w2980 = w2084 ~| w2783;
assign w2981 = ~w2783;
assign w2982 = w2784 & w2785;
assign w2983 = w1551 & w2786;
assign w2984 = w2226 ~| w2787;
assign w2985 = w2713 ~^ w2789;
assign w2986 = ~w2790;
assign w2987 = w2791 & w2792;
assign w2988 = w2790 ~^ w2793;
assign w2989 = ~w2794;
assign w2990 = w2327 & w2795;
assign w2991 = w2332 ^ w2796;
assign w2992 = w2334 ~| w2796;
assign w2993 = w2421 ~^ w2797;
assign w2994 = w2766 | w2798;
assign w2995 = w2338 | w2800;
assign w2996 = w2568 & w2802;
assign w2997 = w2572 ~^ w2806;
assign w2998 = w2572 ~| w2806;
assign w2999 = w2571 | w2807;
assign w3000 = w2734 ^ w2809;
assign w3001 = w2577 | w2810;
assign w3002 = w2809 & w2811;
assign w3003 = w2809 ~| w2811;
assign w3004 = w2580 | w2812;
assign out1[0] = w2464 ~^ w2813;
assign w3005 = w2396 & w2815;
assign w3006 = w2272 ^ w2816;
assign w3007 = w2591 ~^ w2817;
assign w3008 = w2121 | w2819;
assign w3009 = w2586 | w2821;
assign w3010 = w1862 ~^ w2822;
assign w3011 = w1862 | w2824;
assign w3012 = w1873 | w2827;
assign w3013 = w1876 ~^ w2828;
assign w3014 = w2132 ~| w2828;
assign w3015 = ~w2828;
assign w3016 = w2829 & w2830;
assign w3017 = w1567 & w2831;
assign w3018 = w2356 ~| w2832;
assign w3019 = w2513 ~^ w2834;
assign w3020 = w2513 | w2835;
assign w3021 = w2635 | w2836;
assign w3022 = w2789 | w2837;
assign w3023 = w2789 & w2837;
assign w3024 = ~w2838;
assign w3025 = w2839 & w2840;
assign w3026 = w2838 ~^ w2841;
assign w3027 = ~w2842;
assign w3028 = w2374 & w2843;
assign w3029 = w2379 ^ w2844;
assign w3030 = w2381 ~| w2844;
assign w3031 = w2799 ~^ w2845;
assign w3032 = w2799 & w2845;
assign w3033 = w2799 ~| w2845;
assign w3034 = w2385 | w2846;
assign w3035 = w2611 & w2848;
assign w3036 = w2615 ~^ w2852;
assign w3037 = w2615 ~| w2852;
assign w3038 = w2614 | w2853;
assign w3039 = w1208 & w2855;
assign w3040 = w2405 & w2856;
assign w3041 = ~w2857;
assign w3042 = ~w2858;
assign w3043 = w2624 & w2859;
assign w3044 = w2653 ~^ w2861;
assign w3045 = w2653 | w2862;
assign w3046 = w1666 | w2863;
assign w3047 = w1659 ~^ w2864;
assign w3048 = w1909 ~| w2864;
assign w3049 = w1909 & w2864;
assign w3050 = w2634 | w2866;
assign w3051 = w2758 & w2868;
assign w3052 = w2640 & w2869;
assign w3053 = w2640 ~| w2869;
assign w3054 = w2626 ~^ w2870;
assign w3055 = w2627 | w2870;
assign w3056 = w2176 ~^ w2871;
assign w3057 = w2424 ~^ w2873;
assign w3058 = w2424 ~| w2873;
assign w3059 = ~w2873;
assign w3060 = w1201 & w2874;
assign w3061 = w2167 | w2875;
assign w3062 = w2648 ^ w2877;
assign w3063 = w2650 ~| w2877;
assign w3064 = w1280 & w2881;
assign w3065 = w2435 & w2882;
assign w3066 = ~w2883;
assign w3067 = w2658 & w2884;
assign w3068 = w2686 ~^ w2886;
assign w3069 = w2686 | w2887;
assign w3070 = w1708 | w2888;
assign w3071 = w1701 ~^ w2889;
assign w3072 = w1951 ~| w2889;
assign w3073 = w1951 & w2889;
assign w3074 = ~w2890;
assign w3075 = w2668 | w2891;
assign w3076 = w2741 ~| w2892;
assign w3077 = w2673 & w2893;
assign w3078 = w2673 ~| w2893;
assign w3079 = w2660 ~^ w2894;
assign w3080 = w2661 | w2894;
assign w3081 = w2217 ~^ w2895;
assign w3082 = w2454 ~^ w2897;
assign w3083 = w2454 ~| w2897;
assign w3084 = ~w2897;
assign w3085 = w1273 & w2898;
assign w3086 = w2208 | w2899;
assign w3087 = w2092 ~| w2902;
assign w3088 = w2681 ^ w2904;
assign w3089 = w2683 ~| w2904;
assign w3090 = w2816 ~| w2909;
assign w3091 = w2739 ^ w2910;
assign w3092 = w2697 ~| w2910;
assign w3093 = w2697 & w2910;
assign w3094 = w1552 & w2911;
assign w3095 = w2548 & w2912;
assign w3096 = ~w2913;
assign w3097 = w2621 | w2914;
assign w3098 = w2699 ^ w2915;
assign w3099 = w2820 ~| w2915;
assign w3100 = w2820 & w2915;
assign w3101 = w1352 & w2916;
assign w3102 = w2480 & w2917;
assign w3103 = w2521 ~^ w2918;
assign w3104 = ~w2920;
assign w3105 = w2702 & w2921;
assign w3106 = w2733 ~^ w2923;
assign w3107 = w2733 | w2924;
assign w3108 = w1753 | w2925;
assign w3109 = w1746 ~^ w2926;
assign w3110 = w2000 ~| w2926;
assign w3111 = w2000 & w2926;
assign w3112 = w2890 ~| w2927;
assign w3113 = ~w2927;
assign w3114 = w2712 | w2928;
assign w3115 = w2717 & w2929;
assign w3116 = w2717 ~| w2929;
assign w3117 = w2704 ~^ w2930;
assign w3118 = w2705 | w2930;
assign w3119 = w2265 ~^ w2931;
assign w3120 = w2499 ~^ w2933;
assign w3121 = w2499 ~| w2933;
assign w3122 = ~w2933;
assign w3123 = w1345 & w2934;
assign w3124 = w2256 | w2935;
assign w3125 = w2722 | w2937;
assign w3126 = w2767 ~^ w2938;
assign w3127 = w2728 ^ w2940;
assign w3128 = w2730 ~| w2940;
assign w3129 = w1426 & w2945;
assign w3130 = w2518 & w2946;
assign w3131 = w2751 | w2947;
assign w3132 = ~w2947;
assign w3133 = w2669 | w2949;
assign w3134 = ~w2950;
assign w3135 = w2743 & w2951;
assign w3136 = w2776 ~^ w2953;
assign w3137 = w2776 | w2954;
assign w3138 = w1795 | w2955;
assign w3139 = w1788 ~^ w2956;
assign w3140 = w2043 ~| w2956;
assign w3141 = w2043 & w2956;
assign w3142 = w2754 | w2958;
assign w3143 = w2857 ~^ w2959;
assign w3144 = ~w2959;
assign w3145 = w2756 | w2960;
assign w3146 = w2636 ~^ w2961;
assign w3147 = w2762 & w2962;
assign w3148 = w2762 ~| w2962;
assign w3149 = w2745 ~^ w2963;
assign w3150 = w2746 | w2963;
assign w3151 = w2308 ~^ w2964;
assign w3152 = w2538 ~^ w2966;
assign w3153 = w2538 ~| w2966;
assign w3154 = ~w2966;
assign w3155 = w1419 & w2967;
assign w3156 = w2299 | w2968;
assign w3157 = w2644 & w2969;
assign w3158 = w2771 ^ w2972;
assign w3159 = w2773 ~| w2972;
assign w3160 = ~w2976;
assign w3161 = w2778 & w2977;
assign w3162 = w2808 ~^ w2979;
assign w3163 = w2808 | w2980;
assign w3164 = w1831 | w2981;
assign w3165 = w1824 ~^ w2982;
assign w3166 = w2077 ~| w2982;
assign w3167 = w2077 & w2982;
assign w3168 = w2957 ~^ w2983;
assign w3169 = w2865 & w2983;
assign w3170 = w2865 | w2983;
assign w3171 = w2788 | w2984;
assign w3172 = w2837 ~^ w2985;
assign w3173 = w2793 & w2986;
assign w3174 = w2793 ~| w2986;
assign w3175 = w2780 ~^ w2987;
assign w3176 = w2781 | w2987;
assign w3177 = w2342 ~^ w2988;
assign w3178 = w2567 ~^ w2990;
assign w3179 = w2567 ~| w2990;
assign w3180 = ~w2990;
assign w3181 = w1545 & w2991;
assign w3182 = w2333 | w2992;
assign w3183 = w2803 ^ w2996;
assign w3184 = w2805 ~| w2996;
assign w3185 = w2811 ~^ w3000;
assign w3186 = w2944 ^ w3001;
assign w3187 = w2734 ~| w3003;
assign w3188 = w3001 & w3004;
assign w3189 = w3001 ~| w3004;
assign w3190 = w2814 | w3005;
assign w3191 = w2687 ~^ w3006;
assign w3192 = w1568 & w3007;
assign w3193 = w2591 & w3008;
assign w3194 = w2948 ~^ w3009;
assign w3195 = ~w3010;
assign w3196 = w2823 & w3011;
assign w3197 = w2854 ~^ w3013;
assign w3198 = w2854 | w3014;
assign w3199 = w1876 | w3015;
assign w3200 = w1869 ~^ w3016;
assign w3201 = w2125 ~| w3016;
assign w3202 = w2125 & w3016;
assign w3203 = w2927 ~^ w3017;
assign w3204 = ~w3017;
assign w3205 = w2833 | w3018;
assign w3206 = w3020 & w3021;
assign w3207 = w2713 & w3022;
assign w3208 = w2841 & w3024;
assign w3209 = w2841 ~| w3024;
assign w3210 = w2825 ~^ w3025;
assign w3211 = w2826 | w3025;
assign w3212 = w2389 ~^ w3026;
assign w3213 = w2610 ~^ w3028;
assign w3214 = w2610 ~| w3028;
assign w3215 = ~w3028;
assign w3216 = w1561 & w3029;
assign w3217 = w2380 | w3030;
assign w3218 = w2994 ~^ w3031;
assign w3219 = w2994 ~| w3033;
assign w3220 = w2849 ^ w3035;
assign w3221 = w2851 ~| w3035;
assign w3222 = w2619 | w3040;
assign w3223 = ~w3042;
assign w3224 = w2641 ~^ w3043;
assign w3225 = w2872 ~| w3043;
assign w3226 = w2872 & w3043;
assign w3227 = w3045 & w3046;
assign w3228 = w2415 ~^ w3047;
assign w3229 = w2415 ~| w3049;
assign w3230 = w1200 & w3050;
assign w3231 = w2867 | w3051;
assign w3232 = w2176 ~| w3052;
assign w3233 = w2878 ~^ w3054;
assign w3234 = w2880 & w3054;
assign w3235 = w2860 & w3055;
assign w3236 = w1205 & w3056;
assign w3237 = w2876 ~^ w3057;
assign w3238 = w2646 | w3059;
assign w3239 = w1207 & w3061;
assign w3240 = w1881 & w3062;
assign w3241 = w2649 | w3063;
assign w3242 = w2655 | w3065;
assign w3243 = ~w3066;
assign w3244 = w2674 ~^ w3067;
assign w3245 = w2896 ~| w3067;
assign w3246 = w2896 & w3067;
assign w3247 = w3069 & w3070;
assign w3248 = w2445 ~^ w3071;
assign w3249 = w2445 ~| w3073;
assign w3250 = w1272 & w3075;
assign w3251 = w2217 ~| w3077;
assign w3252 = w2905 ~^ w3079;
assign w3253 = w2907 & w3079;
assign w3254 = w2885 & w3080;
assign w3255 = w1277 & w3081;
assign w3256 = w2903 ~^ w3082;
assign w3257 = w2679 | w3084;
assign w3258 = w1279 & w3086;
assign w3259 = w2901 | w3087;
assign w3260 = w1923 & w3088;
assign w3261 = w2682 | w3089;
assign w3262 = w2908 | w3090;
assign w3263 = w2697 ~^ w3091;
assign w3264 = w2739 ~| w3092;
assign w3265 = w2690 | w3095;
assign w3266 = ~w3096;
assign w3267 = w2820 ~^ w3098;
assign w3268 = w2699 ~| w3099;
assign w3269 = w2695 | w3102;
assign w3270 = w2947 ~^ w3103;
assign w3271 = ~w3104;
assign w3272 = w2718 ~^ w3105;
assign w3273 = w2932 ~| w3105;
assign w3274 = w2932 & w3105;
assign w3275 = w3107 & w3108;
assign w3276 = w2490 ~^ w3109;
assign w3277 = w2490 ~| w3111;
assign w3278 = w3074 | w3113;
assign w3279 = w1344 & w3114;
assign w3280 = w2265 ~| w3115;
assign w3281 = w2941 ~^ w3117;
assign w3282 = w2943 & w3117;
assign w3283 = w2922 & w3118;
assign w3284 = w1349 & w3119;
assign w3285 = w2939 ~^ w3120;
assign w3286 = w2726 | w3122;
assign w3287 = w3085 ~^ w3123;
assign w3288 = w3085 | w3123;
assign w3289 = w3085 & w3123;
assign w3290 = w1351 & w3124;
assign w3291 = w2223 ~^ w3125;
assign w3292 = w2900 ~^ w3126;
assign w3293 = ~w3126;
assign w3294 = w1965 & w3127;
assign w3295 = w2729 | w3128;
assign w3296 = w3094 ~^ w3129;
assign w3297 = w3039 | w3129;
assign w3298 = w3039 & w3129;
assign w3299 = w2737 | w3130;
assign w3300 = w2918 & w3131;
assign w3301 = w2521 ~| w3132;
assign w3302 = w3009 & w3133;
assign w3303 = ~w3134;
assign w3304 = w2763 ~^ w3135;
assign w3305 = w2965 ~| w3135;
assign w3306 = w2965 & w3135;
assign w3307 = w3137 & w3138;
assign w3308 = w2529 ~^ w3139;
assign w3309 = w2529 ~| w3141;
assign w3310 = w1418 & w3142;
assign w3311 = w3019 ~^ w3143;
assign w3312 = w3019 | w3144;
assign w3313 = w3019 & w3144;
assign w3314 = w2919 ~^ w3145;
assign w3315 = w2919 & w3145;
assign w3316 = w2919 | w3145;
assign w3317 = ~w3146;
assign w3318 = w2308 ~| w3147;
assign w3319 = w2973 ~^ w3149;
assign w3320 = w2975 & w3149;
assign w3321 = w2952 & w3150;
assign w3322 = w1423 & w3151;
assign w3323 = w2971 ~^ w3152;
assign w3324 = w2769 | w3154;
assign w3325 = ~w3155;
assign w3326 = w1425 & w3156;
assign w3327 = w2970 | w3157;
assign w3328 = w2014 & w3158;
assign w3329 = w2772 | w3159;
assign w3330 = ~w3160;
assign w3331 = w2794 ~^ w3161;
assign w3332 = w2989 ~| w3161;
assign w3333 = w2989 & w3161;
assign w3334 = w3163 & w3164;
assign w3335 = w2558 ~^ w3165;
assign w3336 = w2558 ~| w3167;
assign w3337 = w2865 ~^ w3168;
assign w3338 = w2957 & w3170;
assign w3339 = w1544 & w3171;
assign w3340 = ~w3172;
assign w3341 = w2342 ~| w3173;
assign w3342 = w2997 ~^ w3175;
assign w3343 = w2999 & w3175;
assign w3344 = w2978 & w3176;
assign w3345 = w1549 & w3177;
assign w3346 = w2995 ~^ w3178;
assign w3347 = w2801 | w3180;
assign w3348 = w3155 ~^ w3181;
assign w3349 = ~w3181;
assign w3350 = w1551 & w3182;
assign w3351 = w2091 & w3183;
assign w3352 = w2804 | w3184;
assign w3353 = w3004 ~^ w3186;
assign w3354 = w3002 | w3187;
assign w3355 = w2944 ~| w3189;
assign w3356 = w2508 ~^ w3191;
assign w3357 = w2271 ~| w3191;
assign w3358 = w2271 & w3191;
assign w3359 = w2818 | w3193;
assign w3360 = ~w3194;
assign w3361 = ~w3195;
assign w3362 = w2842 ~^ w3196;
assign w3363 = w3027 ~| w3196;
assign w3364 = w3027 & w3196;
assign w3365 = w3198 & w3199;
assign w3366 = w2601 ~^ w3200;
assign w3367 = w2601 ~| w3202;
assign w3368 = w2890 ~^ w3203;
assign w3369 = w3112 | w3204;
assign w3370 = w1560 & w3205;
assign w3371 = w3146 ~^ w3206;
assign w3372 = w3023 | w3207;
assign w3373 = w2389 ~| w3208;
assign w3374 = w3036 ~^ w3210;
assign w3375 = w3038 & w3210;
assign w3376 = w3012 & w3211;
assign w3377 = w1565 & w3212;
assign w3378 = w3034 ~^ w3213;
assign w3379 = w2847 | w3215;
assign w3380 = w1567 & w3217;
assign w3381 = ~w3218;
assign w3382 = w3032 | w3219;
assign w3383 = w2095 & w3220;
assign w3384 = w2850 | w3221;
assign w3385 = w1200 & w3222;
assign w3386 = w3224 ~^ w3227;
assign w3387 = w3226 ~| w3227;
assign w3388 = w1208 & w3228;
assign w3389 = w3048 | w3229;
assign w3390 = w3053 | w3232;
assign w3391 = w1211 & w3233;
assign w3392 = w2879 | w3234;
assign w3393 = w2858 ~^ w3235;
assign w3394 = w3223 ~| w3235;
assign w3395 = ~w3235;
assign w3396 = w1209 & w3237;
assign w3397 = w2876 & w3238;
assign w3398 = w1209 & w3241;
assign w3399 = w1272 & w3242;
assign w3400 = w3244 ~^ w3247;
assign w3401 = w3246 ~| w3247;
assign w3402 = w1280 & w3248;
assign w3403 = w3072 | w3249;
assign w3404 = w3230 ~^ w3250;
assign w3405 = w3078 | w3251;
assign w3406 = w1283 & w3252;
assign w3407 = w2906 | w3253;
assign w3408 = w2883 ~^ w3254;
assign w3409 = w3243 ~| w3254;
assign w3410 = ~w3254;
assign w3411 = w1281 & w3256;
assign w3412 = w2903 & w3257;
assign w3413 = w2993 ~^ w3258;
assign w3414 = w2421 ~| w3258;
assign w3415 = w2421 & w3258;
assign w3416 = w2578 ~^ w3259;
assign w3417 = w1281 & w3261;
assign w3418 = w3096 ~^ w3263;
assign w3419 = ~w3263;
assign w3420 = w3093 | w3264;
assign w3421 = w1544 & w3265;
assign w3422 = w3263 | w3266;
assign w3423 = w3097 ^ w3267;
assign w3424 = ~w3267;
assign w3425 = w3100 | w3268;
assign w3426 = w1344 & w3269;
assign w3427 = ~w3270;
assign w3428 = w3272 ~^ w3275;
assign w3429 = w3274 ~| w3275;
assign w3430 = w1352 & w3276;
assign w3431 = w3110 | w3277;
assign w3432 = w3064 ~^ w3279;
assign w3433 = w3101 | w3279;
assign w3434 = w3101 & w3279;
assign w3435 = w3116 | w3280;
assign w3436 = w1355 & w3281;
assign w3437 = w2942 | w3282;
assign w3438 = w2920 ~^ w3283;
assign w3439 = w3271 ~| w3283;
assign w3440 = ~w3283;
assign w3441 = w1353 & w3285;
assign w3442 = w2939 & w3286;
assign w3443 = w3216 ~^ w3287;
assign w3444 = w3216 & w3288;
assign w3445 = w3239 ~^ w3290;
assign w3446 = w3239 | w3290;
assign w3447 = w3239 & w3290;
assign w3448 = w3218 ~^ w3292;
assign w3449 = w3218 & w3293;
assign w3450 = w1353 & w3295;
assign w3451 = w3039 ~^ w3296;
assign w3452 = w3094 & w3297;
assign w3453 = w1418 & w3299;
assign w3454 = w3300 | w3301;
assign w3455 = w3076 | w3302;
assign w3456 = w3304 ~^ w3307;
assign w3457 = w3306 ~| w3307;
assign w3458 = w1426 & w3308;
assign w3459 = w3140 | w3309;
assign w3460 = w3310 ~^ in5[5];
assign w3461 = w3041 | w3313;
assign w3462 = ~w3317;
assign w3463 = w3148 | w3318;
assign w3464 = w1429 & w3319;
assign w3465 = w2974 | w3320;
assign w3466 = w2950 ~^ w3321;
assign w3467 = w3303 ~| w3321;
assign w3468 = ~w3321;
assign w3469 = w3236 ~^ w3322;
assign w3470 = w1427 & w3323;
assign w3471 = w2971 & w3324;
assign w3472 = ~w3328;
assign w3473 = w1427 & w3329;
assign w3474 = w3331 ~^ w3334;
assign w3475 = w3333 ~| w3334;
assign w3476 = w1552 & w3335;
assign w3477 = w3166 | w3336;
assign w3478 = w3314 ~^ w3337;
assign w3479 = w3316 & w3337;
assign w3480 = w3169 | w3338;
assign w3481 = w3230 | w3339;
assign w3482 = w3230 & w3339;
assign w3483 = w3194 ~| w3340;
assign w3484 = w3174 | w3341;
assign w3485 = w1555 & w3342;
assign w3486 = w2998 | w3343;
assign w3487 = w2976 ~^ w3344;
assign w3488 = w3330 ~| w3344;
assign w3489 = ~w3344;
assign w3490 = w3236 | w3345;
assign w3491 = w3236 & w3345;
assign w3492 = w1553 & w3346;
assign w3493 = w2995 & w3347;
assign w3494 = w3325 | w3349;
assign w3495 = w1553 & w3352;
assign w3496 = w3353 ~^ w3354;
assign w3497 = w3353 & w3354;
assign w3498 = w3353 | w3354;
assign w3499 = w3188 | w3355;
assign w3500 = w3185 ~^ w3356;
assign w3501 = w3185 & w3356;
assign w3502 = w3185 | w3356;
assign w3503 = w2397 ~| w3357;
assign w3504 = w1560 & w3359;
assign w3505 = w3172 | w3360;
assign w3506 = w3362 ~^ w3365;
assign w3507 = w3364 ~| w3365;
assign w3508 = w1568 & w3366;
assign w3509 = w3201 | w3367;
assign w3510 = ~w3368;
assign w3511 = w3278 & w3369;
assign w3512 = in5[5] | w3370;
assign w3513 = in5[5] & w3370;
assign w3514 = w3368 ~^ w3371;
assign w3515 = ~w3372;
assign w3516 = w3209 | w3373;
assign w3517 = w1571 & w3374;
assign w3518 = w3037 | w3375;
assign w3519 = w3010 ~^ w3376;
assign w3520 = w3361 ~| w3376;
assign w3521 = ~w3376;
assign w3522 = ~w3377;
assign w3523 = w1569 & w3378;
assign w3524 = w3034 & w3379;
assign w3525 = w3350 ~^ w3380;
assign w3526 = w3350 & w3380;
assign w3527 = w3350 ~| w3380;
assign w3528 = w3126 & w3381;
assign w3529 = w3327 ~^ w3382;
assign w3530 = w1569 & w3384;
assign w3531 = in5[6] | w3385;
assign w3532 = in5[6] & w3385;
assign w3533 = w1206 & w3386;
assign w3534 = w3225 | w3387;
assign w3535 = w1197 & w3389;
assign w3536 = w1203 & w3390;
assign w3537 = w1202 & w3392;
assign w3538 = w3044 ~^ w3393;
assign w3539 = w3042 | w3395;
assign w3540 = w3058 | w3397;
assign w3541 = w1278 & w3400;
assign w3542 = w3245 | w3401;
assign w3543 = w1269 & w3403;
assign w3544 = w3339 ~^ w3404;
assign w3545 = w1275 & w3405;
assign w3546 = ~w3406;
assign w3547 = w1274 & w3407;
assign w3548 = w3068 ~^ w3408;
assign w3549 = w3066 | w3410;
assign w3550 = w3396 & w3411;
assign w3551 = w3396 | w3411;
assign w3552 = w3083 | w3412;
assign w3553 = w2797 ~| w3414;
assign w3554 = w2574 ~^ w3416;
assign w3555 = w3060 ~^ w3417;
assign w3556 = w3060 & w3417;
assign w3557 = w3060 | w3417;
assign w3558 = w3096 ~| w3419;
assign w3559 = ~w3420;
assign w3560 = w3311 ~^ w3423;
assign w3561 = w3311 & w3424;
assign w3562 = w3311 ~| w3424;
assign w3563 = ~w3425;
assign w3564 = w3421 ~^ w3426;
assign w3565 = w1350 & w3428;
assign w3566 = w3273 | w3429;
assign w3567 = w3402 & w3430;
assign w3568 = w3402 | w3430;
assign w3569 = w1341 & w3431;
assign w3570 = w3101 ~^ w3432;
assign w3571 = w3064 & w3433;
assign w3572 = w1347 & w3435;
assign w3573 = ~w3436;
assign w3574 = w1346 & w3437;
assign w3575 = w3106 ~^ w3438;
assign w3576 = w3104 | w3440;
assign w3577 = w3411 ~^ w3441;
assign w3578 = w3121 | w3442;
assign w3579 = w3289 | w3444;
assign w3580 = w3326 ~^ w3445;
assign w3581 = w3326 & w3446;
assign w3582 = w2900 ~| w3449;
assign w3583 = ~w3451;
assign w3584 = w3298 | w3452;
assign w3585 = w3453 ~^ in5[6];
assign w3586 = w3172 ~^ w3454;
assign w3587 = w1424 & w3456;
assign w3588 = w3305 | w3457;
assign w3589 = w1415 & w3459;
assign w3590 = w3370 ~^ w3460;
assign w3591 = w3312 & w3461;
assign w3592 = w3368 ~| w3462;
assign w3593 = w1421 & w3463;
assign w3594 = w1420 & w3465;
assign w3595 = w3136 ~^ w3466;
assign w3596 = w3134 | w3468;
assign w3597 = w3345 ~^ w3469;
assign w3598 = ~w3470;
assign w3599 = w3153 | w3471;
assign w3600 = w3398 ~^ w3473;
assign w3601 = w3398 & w3473;
assign w3602 = w3398 | w3473;
assign w3603 = w1550 & w3474;
assign w3604 = w3332 | w3475;
assign w3605 = w3458 ~^ w3476;
assign w3606 = w3388 & w3476;
assign w3607 = w3388 | w3476;
assign w3608 = w1541 & w3477;
assign w3609 = w3425 ~| w3478;
assign w3610 = ~w3478;
assign w3611 = w3315 | w3479;
assign w3612 = w3192 ~^ w3480;
assign w3613 = w3192 & w3480;
assign w3614 = w3192 | w3480;
assign w3615 = w3250 & w3481;
assign w3616 = w1547 & w3484;
assign w3617 = w1546 & w3486;
assign w3618 = w3162 ~^ w3487;
assign w3619 = w3160 | w3489;
assign w3620 = w3322 & w3490;
assign w3621 = ~w3492;
assign w3622 = w3179 | w3493;
assign w3623 = w3262 ~^ w3496;
assign w3624 = w3262 & w3498;
assign w3625 = w3270 ~^ w3499;
assign w3626 = w3427 ~| w3499;
assign w3627 = ~w3499;
assign out1[1] = w3190 ~^ w3500;
assign w3628 = w3190 & w3502;
assign w3629 = w3358 | w3503;
assign w3630 = w3421 & w3504;
assign w3631 = w3421 | w3504;
assign w3632 = w3454 & w3505;
assign w3633 = w1566 & w3506;
assign w3634 = w3363 | w3507;
assign w3635 = w3430 ~^ w3508;
assign w3636 = w1557 & w3509;
assign w3637 = w3317 | w3510;
assign w3638 = w3310 & w3512;
assign w3639 = w3511 ~^ w3515;
assign w3640 = w1563 & w3516;
assign w3641 = ~w3517;
assign w3642 = w1562 & w3518;
assign w3643 = w3197 ~^ w3519;
assign w3644 = w3195 | w3521;
assign w3645 = w3492 ~^ w3523;
assign w3646 = ~w3523;
assign w3647 = w3214 | w3524;
assign w3648 = w3494 ~^ w3525;
assign w3649 = w3494 ~| w3527;
assign w3650 = ~w3529;
assign w3651 = w3348 ~^ w3530;
assign w3652 = ~w3530;
assign w3653 = w3453 & w3531;
assign w3654 = ~w3533;
assign w3655 = w1201 & w3534;
assign w3656 = w3255 ~^ w3535;
assign w3657 = w3284 | w3535;
assign w3658 = w3284 & w3535;
assign w3659 = w3485 & w3536;
assign w3660 = w3485 | w3536;
assign w3661 = ~w3537;
assign w3662 = w1210 & w3538;
assign w3663 = w3044 & w3539;
assign w3664 = w1882 & w3540;
assign w3665 = w3533 ~| w3541;
assign w3666 = ~w3541;
assign w3667 = w1273 & w3542;
assign w3668 = w3372 ~| w3544;
assign w3669 = ~w3544;
assign w3670 = w3391 ~^ w3545;
assign w3671 = w3464 & w3545;
assign w3672 = w3464 | w3545;
assign w3673 = w1282 & w3548;
assign w3674 = w3068 & w3549;
assign w3675 = w3441 & w3551;
assign w3676 = w1924 & w3552;
assign w3677 = w3415 | w3553;
assign w3678 = w3450 ~^ w3555;
assign w3679 = w3450 & w3557;
assign w3680 = w3097 ~| w3561;
assign w3681 = w3504 ^ w3564;
assign w3682 = w3541 ~^ w3565;
assign w3683 = ~w3565;
assign w3684 = w1345 & w3566;
assign w3685 = w3508 & w3568;
assign w3686 = w3543 ~^ w3569;
assign w3687 = ~w3570;
assign w3688 = w3434 | w3571;
assign w3689 = w3406 ~^ w3572;
assign w3690 = ~w3572;
assign w3691 = w1354 & w3575;
assign w3692 = w3106 & w3576;
assign w3693 = w3396 ~^ w3577;
assign w3694 = w1967 & w3578;
assign w3695 = w2936 ~^ w3579;
assign w3696 = w2936 & w3579;
assign w3697 = w2936 | w3579;
assign w3698 = ~w3580;
assign w3699 = w3447 | w3581;
assign w3700 = w3528 ~| w3582;
assign w3701 = w3385 ~^ w3585;
assign w3702 = w3194 ~^ w3586;
assign w3703 = w1419 & w3588;
assign w3704 = ~w3589;
assign w3705 = w3451 ~^ w3590;
assign w3706 = w3451 ~| w3590;
assign w3707 = ~w3590;
assign w3708 = w3425 ~^ w3591;
assign w3709 = w3206 | w3592;
assign w3710 = w3517 ~^ w3593;
assign w3711 = ~w3593;
assign w3712 = ~w3594;
assign w3713 = w1428 & w3595;
assign w3714 = w3136 & w3596;
assign w3715 = ~w3597;
assign w3716 = w2016 & w3599;
assign w3717 = w3495 ~^ w3600;
assign w3718 = w3495 & w3602;
assign w3719 = ~w3603;
assign w3720 = w1545 & w3604;
assign w3721 = w3388 ~^ w3605;
assign w3722 = w3458 & w3607;
assign w3723 = w3589 ~^ w3608;
assign w3724 = ~w3608;
assign w3725 = w3591 | w3609;
assign w3726 = w3563 | w3610;
assign w3727 = w3455 & w3611;
assign w3728 = w3455 ~| w3611;
assign w3729 = w3231 ~^ w3612;
assign w3730 = w3231 & w3614;
assign w3731 = w3482 | w3615;
assign w3732 = w3485 ~^ w3616;
assign w3733 = ~w3617;
assign w3734 = w1554 & w3618;
assign w3735 = w3162 & w3619;
assign w3736 = w3491 | w3620;
assign w3737 = w2094 & w3622;
assign w3738 = ~w3623;
assign w3739 = w3497 | w3624;
assign w3740 = w3420 ~^ w3625;
assign w3741 = w3559 | w3626;
assign w3742 = w3270 | w3627;
assign w3743 = w3501 | w3628;
assign w3744 = w3418 ~^ w3629;
assign w3745 = w3422 & w3629;
assign w3746 = w3426 & w3631;
assign w3747 = w3483 | w3632;
assign w3748 = w3603 ~^ w3633;
assign w3749 = ~w3633;
assign w3750 = w1561 & w3634;
assign w3751 = w3402 ~^ w3635;
assign w3752 = w3543 & w3636;
assign w3753 = w3543 | w3636;
assign w3754 = w3513 | w3638;
assign w3755 = w3544 ~^ w3639;
assign w3756 = w3406 ~| w3640;
assign w3757 = ~w3640;
assign w3758 = w1570 & w3643;
assign w3759 = w3197 & w3644;
assign w3760 = w3621 | w3646;
assign w3761 = w2098 & w3647;
assign w3762 = ~w3648;
assign w3763 = w3526 | w3649;
assign w3764 = w3532 | w3653;
assign w3765 = w3284 ~^ w3656;
assign w3766 = w3255 & w3657;
assign w3767 = w3616 & w3660;
assign w3768 = w3547 ~^ w3662;
assign w3769 = w3394 | w3663;
assign w3770 = w3260 ~^ w3664;
assign w3771 = w3260 | w3664;
assign w3772 = w3260 & w3664;
assign w3773 = w3654 | w3666;
assign w3774 = w3655 & w3667;
assign w3775 = w3655 | w3667;
assign w3776 = w3511 | w3668;
assign w3777 = w3515 | w3669;
assign w3778 = w3464 ^ w3670;
assign w3779 = w3391 & w3672;
assign w3780 = w3574 ~^ w3673;
assign w3781 = w3642 | w3673;
assign w3782 = w3642 & w3673;
assign w3783 = w3409 | w3674;
assign w3784 = w3550 | w3675;
assign w3785 = w3294 ~^ w3676;
assign w3786 = w3294 | w3676;
assign w3787 = w3294 & w3676;
assign w3788 = w3556 | w3679;
assign w3789 = w3562 | w3680;
assign w3790 = w3533 ~^ w3682;
assign w3791 = w3665 | w3683;
assign w3792 = w3645 ~^ w3684;
assign w3793 = ~w3684;
assign w3794 = w3567 | w3685;
assign w3795 = w3636 ~^ w3686;
assign w3796 = w3584 ~^ w3688;
assign w3797 = w3584 | w3688;
assign w3798 = w3584 & w3688;
assign w3799 = w3640 ~^ w3689;
assign w3800 = ~w3691;
assign w3801 = w3439 | w3692;
assign w3802 = ~w3694;
assign w3803 = w3291 ~^ w3699;
assign w3804 = w3125 | w3699;
assign w3805 = w3125 & w3699;
assign w3806 = w3554 ~^ w3700;
assign w3807 = w3681 ^ w3701;
assign w3808 = w3514 | w3702;
assign w3809 = w3514 & w3702;
assign w3810 = w3470 ~^ w3703;
assign w3811 = ~w3703;
assign w3812 = w3570 ~^ w3705;
assign w3813 = w3687 | w3706;
assign w3814 = w3583 | w3707;
assign w3815 = w3478 ~^ w3708;
assign w3816 = w3637 & w3709;
assign w3817 = w3641 | w3711;
assign w3818 = w3547 | w3713;
assign w3819 = w3547 & w3713;
assign w3820 = w3467 | w3714;
assign w3821 = ~w3717;
assign w3822 = w3601 | w3718;
assign w3823 = w3470 ~| w3720;
assign w3824 = ~w3720;
assign w3825 = w3606 | w3722;
assign w3826 = w3377 ~^ w3723;
assign w3827 = w3522 ~| w3723;
assign w3828 = ~w3723;
assign w3829 = w3704 | w3724;
assign w3830 = w3725 & w3726;
assign w3831 = w3613 | w3730;
assign w3832 = w3399 ~^ w3731;
assign w3833 = ~w3731;
assign w3834 = w3536 ~^ w3732;
assign w3835 = w3617 ~^ w3734;
assign w3836 = w3537 ~| w3734;
assign w3837 = ~w3734;
assign w3838 = w3488 | w3735;
assign w3839 = ~w3736;
assign w3840 = w3351 ~^ w3737;
assign w3841 = w3240 | w3737;
assign w3842 = w3240 & w3737;
assign w3843 = ~w3739;
assign w3844 = w3739 ~^ w3740;
assign w3845 = w3741 & w3742;
assign w3846 = w3623 ~^ w3744;
assign w3847 = w3738 ~| w3744;
assign w3848 = ~w3744;
assign w3849 = w3558 | w3745;
assign w3850 = w3630 | w3746;
assign w3851 = w3719 | w3749;
assign w3852 = w3667 ~^ w3750;
assign w3853 = w3701 & w3751;
assign w3854 = w3701 ~| w3751;
assign w3855 = w3569 & w3753;
assign w3856 = w3399 ~| w3754;
assign w3857 = w3399 & w3754;
assign w3858 = w3729 ~^ w3755;
assign w3859 = w3729 & w3755;
assign w3860 = w3729 | w3755;
assign w3861 = w3690 | w3756;
assign w3862 = w3546 | w3757;
assign w3863 = w3594 ~^ w3758;
assign w3864 = ~w3758;
assign w3865 = w3520 | w3759;
assign w3866 = w3328 ~^ w3761;
assign w3867 = ~w3761;
assign w3868 = w3677 ~^ w3763;
assign w3869 = w3677 | w3763;
assign w3870 = w3677 & w3763;
assign w3871 = ~w3765;
assign w3872 = w3658 | w3766;
assign w3873 = w3659 | w3767;
assign w3874 = w3713 ~^ w3768;
assign w3875 = w1198 & w3769;
assign w3876 = w3716 ~^ w3770;
assign w3877 = w3716 & w3771;
assign w3878 = w3750 & w3775;
assign w3879 = w3776 & w3777;
assign w3880 = w3671 | w3779;
assign w3881 = w3642 ~^ w3780;
assign w3882 = w3574 & w3781;
assign w3883 = w1270 & w3783;
assign w3884 = ~w3784;
assign w3885 = w3383 ~^ w3785;
assign w3886 = w3383 & w3786;
assign w3887 = w3580 ~^ w3788;
assign w3888 = w3580 ~| w3788;
assign w3889 = ~w3788;
assign w3890 = ~w3789;
assign w3891 = ~w3790;
assign w3892 = w3773 & w3791;
assign w3893 = w3597 ~^ w3795;
assign w3894 = w3597 ~| w3795;
assign w3895 = ~w3795;
assign w3896 = w3721 ~^ w3796;
assign w3897 = w3721 & w3797;
assign w3898 = w1342 & w3801;
assign w3899 = w3760 ~| w3802;
assign w3900 = w3760 & w3802;
assign w3901 = w2223 & w3804;
assign w3902 = w3751 ~^ w3807;
assign w3903 = w3720 ~^ w3810;
assign w3904 = ~w3812;
assign w3905 = w3813 & w3814;
assign w3906 = w3789 ~^ w3815;
assign w3907 = w3455 ~^ w3816;
assign w3908 = w3728 ~| w3816;
assign w3909 = w3662 & w3818;
assign w3910 = w1416 & w3820;
assign w3911 = w3695 ~^ w3822;
assign w3912 = w3697 & w3822;
assign w3913 = w3811 | w3823;
assign w3914 = w3598 | w3824;
assign w3915 = w3764 ~^ w3826;
assign w3916 = w3377 | w3828;
assign w3917 = w3436 ~^ w3829;
assign w3918 = w3573 | w3829;
assign w3919 = ~w3829;
assign w3920 = w3754 ~^ w3832;
assign w3921 = w3778 ^ w3834;
assign w3922 = w3799 ~| w3834;
assign w3923 = w3799 & w3834;
assign w3924 = w3537 ^ w3835;
assign w3925 = w3733 | w3836;
assign w3926 = w3661 | w3837;
assign w3927 = w1542 & w3838;
assign w3928 = w3240 ~^ w3840;
assign w3929 = w3351 & w3841;
assign w3930 = w3740 ~| w3843;
assign w3931 = w3740 & w3843;
assign w3932 = w3560 ~^ w3844;
assign w3933 = w3809 | w3845;
assign w3934 = w3514 ~^ w3845;
assign out1[2] = w3743 ^ w3846;
assign w3935 = w3623 | w3848;
assign w3936 = w3794 ~^ w3850;
assign w3937 = w3794 & w3850;
assign w3938 = w3794 | w3850;
assign w3939 = w3792 ~^ w3851;
assign w3940 = w3793 ~| w3851;
assign w3941 = w3793 & w3851;
assign w3942 = w3655 ~^ w3852;
assign w3943 = w3681 ~| w3854;
assign w3944 = w3752 | w3855;
assign w3945 = w3833 ~| w3856;
assign w3946 = w3747 ~^ w3858;
assign w3947 = w3747 & w3860;
assign w3948 = w3861 & w3862;
assign w3949 = w3691 ~^ w3863;
assign w3950 = w3800 | w3863;
assign w3951 = ~w3863;
assign w3952 = w3712 | w3864;
assign w3953 = w1558 & w3865;
assign w3954 = w3694 ~^ w3866;
assign w3955 = w3472 | w3867;
assign w3956 = w3803 ~^ w3868;
assign w3957 = w3803 & w3869;
assign w3958 = ~w3872;
assign w3959 = ~w3873;
assign w3960 = w3772 | w3877;
assign w3961 = w3774 | w3878;
assign w3962 = w3831 ^ w3879;
assign w3963 = w3873 ~| w3880;
assign w3964 = ~w3880;
assign w3965 = w3874 & w3881;
assign w3966 = w3874 ~| w3881;
assign w3967 = w3782 | w3882;
assign w3968 = w3875 & w3883;
assign w3969 = w3875 | w3883;
assign w3970 = w3876 ~^ w3885;
assign w3971 = w3876 & w3885;
assign w3972 = w3876 | w3885;
assign w3973 = w3787 | w3886;
assign w3974 = w3413 ~^ w3887;
assign w3975 = w3413 | w3888;
assign w3976 = w3698 | w3889;
assign w3977 = w3815 ~| w3890;
assign w3978 = w3815 & w3890;
assign w3979 = w3715 | w3895;
assign w3980 = w3798 | w3897;
assign w3981 = w3748 ~^ w3898;
assign w3982 = ~w3898;
assign w3983 = w3866 ~| w3900;
assign w3984 = w3805 | w3901;
assign w3985 = w3896 & w3902;
assign w3986 = w3896 ~| w3902;
assign w3987 = w3830 ~^ w3904;
assign w3988 = w3896 ^ w3905;
assign w3989 = w3611 ~^ w3907;
assign w3990 = w3727 | w3908;
assign w3991 = w3819 | w3909;
assign w3992 = w3587 ~^ w3910;
assign w3993 = ~w3911;
assign w3994 = w3696 | w3912;
assign w3995 = w3913 & w3914;
assign w3996 = w3765 ~^ w3915;
assign w3997 = w3871 ~| w3915;
assign w3998 = ~w3915;
assign w3999 = w3764 & w3916;
assign w4000 = w3710 ~^ w3917;
assign w4001 = w3436 ~| w3919;
assign w4002 = w3831 & w3920;
assign w4003 = w3831 ~| w3920;
assign w4004 = w3799 ~^ w3921;
assign w4005 = w3778 ~| w3922;
assign w4006 = w3874 ^ w3924;
assign w4007 = w3925 & w3926;
assign w4008 = w3587 | w3927;
assign w4009 = w3587 & w3927;
assign w4010 = w3784 ~| w3928;
assign w4011 = ~w3928;
assign w4012 = w3842 | w3929;
assign w4013 = w3560 ~| w3931;
assign w4014 = w3849 ~^ w3932;
assign w4015 = w3849 & w3932;
assign w4016 = w3849 | w3932;
assign w4017 = w3808 & w3933;
assign w4018 = w3702 ~^ w3934;
assign w4019 = w3743 & w3935;
assign w4020 = w3825 ~^ w3936;
assign w4021 = w3825 & w3938;
assign w4022 = w3903 ~^ w3939;
assign w4023 = w3903 | w3939;
assign w4024 = w3903 & w3939;
assign w4025 = w3645 ~| w3941;
assign w4026 = ~w3942;
assign w4027 = w3853 | w3943;
assign w4028 = w3872 ~^ w3944;
assign w4029 = w3872 ~| w3944;
assign w4030 = ~w3944;
assign w4031 = w3857 | w3945;
assign w4032 = w3812 ~| w3946;
assign w4033 = ~w3946;
assign w4034 = w3859 | w3947;
assign w4035 = w3880 ^ w3948;
assign w4036 = w3817 ~^ w3949;
assign w4037 = w3691 ~| w3951;
assign w4038 = ~w3952;
assign w4039 = w3883 ~^ w3953;
assign w4040 = w3760 ~^ w3954;
assign w4041 = w3651 ~^ w3955;
assign w4042 = w3652 ~| w3955;
assign w4043 = w3652 & w3955;
assign w4044 = w3870 | w3957;
assign w4045 = w3717 ~^ w3960;
assign w4046 = w3678 & w3960;
assign w4047 = w3678 ~| w3960;
assign w4048 = w3920 ~^ w3962;
assign w4049 = w3948 | w3963;
assign w4050 = w3959 | w3964;
assign w4051 = w3924 ~| w3966;
assign w4052 = w3953 & w3969;
assign w4053 = w3961 ~^ w3970;
assign w4054 = w3961 & w3972;
assign w4055 = w3443 ~^ w3973;
assign w4056 = ~w3974;
assign w4057 = w3975 & w3976;
assign w4058 = w3952 ~^ w3981;
assign w4059 = w3952 | w3982;
assign w4060 = w3899 | w3983;
assign w4061 = w3806 ~^ w3984;
assign w4062 = w3905 ~| w3986;
assign w4063 = w3946 ~^ w3987;
assign w4064 = w3902 ^ w3988;
assign w4065 = ~w3989;
assign w4066 = ~w3990;
assign w4067 = w3967 ~| w3991;
assign w4068 = w3967 & w3991;
assign w4069 = w3927 ~^ w3992;
assign w4070 = w3448 ~^ w3994;
assign w4071 = w3884 ~^ w3995;
assign w4072 = w3765 | w3998;
assign w4073 = w3827 | w3999;
assign w4074 = w3710 | w4001;
assign w4075 = w3879 ~| w4003;
assign w4076 = w3923 | w4005;
assign w4077 = w3881 ~^ w4006;
assign w4078 = w3967 ^ w4007;
assign w4079 = w3910 & w4008;
assign w4080 = w3995 | w4010;
assign w4081 = w3884 | w4011;
assign w4082 = w3973 | w4012;
assign w4083 = w3973 & w4012;
assign w4084 = w3930 | w4013;
assign w4085 = w3989 ~^ w4017;
assign w4086 = w3906 ~^ w4018;
assign w4087 = w3978 ~| w4018;
assign w4088 = w3847 | w4019;
assign w4089 = w3980 ~^ w4020;
assign w4090 = w3980 | w4020;
assign w4091 = w3980 & w4020;
assign w4092 = w3937 | w4021;
assign w4093 = w3940 | w4025;
assign w4094 = w3996 ~^ w4027;
assign w4095 = w3736 ~^ w4028;
assign w4096 = w3839 | w4029;
assign w4097 = w3958 | w4030;
assign w4098 = w3893 ~^ w4031;
assign w4099 = ~w4031;
assign w4100 = w3830 | w4032;
assign w4101 = w3904 | w4033;
assign w4102 = w3873 ~^ w4035;
assign w4103 = ~w4036;
assign w4104 = w3817 | w4037;
assign w4105 = w3898 ~| w4038;
assign w4106 = w3875 ~^ w4039;
assign w4107 = ~w4040;
assign w4108 = ~w4041;
assign w4109 = w3348 ~| w4043;
assign w4110 = w3650 ~^ w4044;
assign w4111 = w3678 ~^ w4045;
assign w4112 = w3821 ~| w4047;
assign w4113 = w3990 | w4048;
assign w4114 = ~w4048;
assign w4115 = w4049 & w4050;
assign w4116 = w3965 | w4051;
assign w4117 = w3968 | w4052;
assign w4118 = w3971 | w4054;
assign w4119 = w4012 ~^ w4055;
assign w4120 = ~w4057;
assign w4121 = w4041 ~^ w4060;
assign w4122 = w4041 ~| w4060;
assign w4123 = ~w4060;
assign w4124 = w3985 | w4062;
assign w4125 = w4063 & w4065;
assign w4126 = w4063 ~| w4065;
assign w4127 = w4048 ~^ w4066;
assign w4128 = w4007 ~| w4067;
assign w4129 = w4058 & w4069;
assign w4130 = w4058 ~| w4069;
assign w4131 = w4057 ~^ w4070;
assign w4132 = w3928 ~^ w4071;
assign w4133 = w4027 & w4072;
assign w4134 = w4000 | w4073;
assign w4135 = w4000 & w4073;
assign w4136 = w3918 & w4074;
assign w4137 = w4002 | w4075;
assign w4138 = w3991 ~^ w4078;
assign w4139 = w4009 | w4079;
assign w4140 = w4080 & w4081;
assign w4141 = w3443 & w4082;
assign w4142 = w4063 ~^ w4085;
assign w4143 = w4084 ~^ w4086;
assign w4144 = w4084 & w4086;
assign w4145 = w4084 | w4086;
assign w4146 = w3977 | w4087;
assign out1[3] = w4014 ~^ w4088;
assign w4147 = w4016 & w4088;
assign w4148 = w4073 ~^ w4092;
assign w4149 = w4040 | w4093;
assign w4150 = ~w4093;
assign w4151 = ~w4094;
assign w4152 = w4004 & w4095;
assign w4153 = w4004 ~| w4095;
assign w4154 = w4096 & w4097;
assign w4155 = w4094 ~^ w4098;
assign w4156 = ~w4098;
assign w4157 = w3894 | w4099;
assign w4158 = w4100 & w4101;
assign w4159 = w4076 ~^ w4102;
assign w4160 = w4076 | w4102;
assign w4161 = w4076 & w4102;
assign w4162 = w3950 & w4104;
assign w4163 = w3748 | w4105;
assign w4164 = w3790 ~^ w4106;
assign w4165 = w3790 ~| w4106;
assign w4166 = ~w4106;
assign w4167 = w4042 | w4109;
assign w4168 = w4046 | w4112;
assign w4169 = w4034 & w4113;
assign w4170 = w4066 ~| w4114;
assign w4171 = w4069 ^ w4115;
assign w4172 = ~w4116;
assign w4173 = w3693 ~| w4117;
assign w4174 = w3693 & w4117;
assign w4175 = w3892 ^ w4117;
assign w4176 = ~w4118;
assign w4177 = w4111 & w4119;
assign w4178 = w4111 ~| w4119;
assign w4179 = w3994 | w4120;
assign w4180 = w3994 & w4120;
assign w4181 = w4118 ~^ w4121;
assign w4182 = w4108 | w4123;
assign w4183 = ~w4124;
assign w4184 = w4017 ~| w4126;
assign w4185 = w4034 ~^ w4127;
assign w4186 = w4068 | w4128;
assign w4187 = w4115 ~| w4130;
assign w4188 = w4053 & w4132;
assign w4189 = w4053 ~| w4132;
assign w4190 = w3997 | w4133;
assign w4191 = w4092 & w4134;
assign w4192 = w4103 & w4136;
assign w4193 = w4103 ~| w4136;
assign w4194 = w4089 ~^ w4137;
assign w4195 = w4090 & w4137;
assign w4196 = w4116 ~^ w4138;
assign w4197 = w4116 ~| w4138;
assign w4198 = ~w4138;
assign w4199 = w3942 ~^ w4139;
assign w4200 = w3942 ~| w4139;
assign w4201 = ~w4139;
assign w4202 = w4119 ^ w4140;
assign w4203 = w4083 | w4141;
assign w4204 = w4142 ~^ w4146;
assign w4205 = w4142 & w4146;
assign w4206 = w4142 | w4146;
assign w4207 = w4015 | w4147;
assign w4208 = w4000 ~^ w4148;
assign w4209 = w4040 ~^ w4150;
assign w4210 = w4107 ~| w4150;
assign w4211 = w4098 ~| w4151;
assign w4212 = w4136 ~^ w4154;
assign w4213 = w4124 ~^ w4155;
assign w4214 = w4094 | w4156;
assign w4215 = w3979 & w4157;
assign w4216 = w4064 ^ w4158;
assign w4217 = w4059 & w4163;
assign w4218 = w4162 ^ w4164;
assign w4219 = w4162 | w4165;
assign w4220 = w3891 | w4166;
assign w4221 = w3648 ~^ w4167;
assign w4222 = w3762 ~| w4167;
assign w4223 = ~w4167;
assign w4224 = w4056 | w4168;
assign w4225 = ~w4168;
assign w4226 = w4169 | w4170;
assign w4227 = w4058 ~^ w4171;
assign w4228 = w3892 ~| w4173;
assign w4229 = w3693 ^ w4175;
assign w4230 = w4122 | w4176;
assign w4231 = w4140 ~| w4178;
assign w4232 = w3448 & w4179;
assign w4233 = ~w4181;
assign w4234 = w4125 | w4184;
assign w4235 = w4064 | w4185;
assign w4236 = w4064 & w4185;
assign w4237 = w4022 ~^ w4186;
assign w4238 = w4023 & w4186;
assign w4239 = w4129 | w4187;
assign w4240 = w4135 | w4191;
assign w4241 = w4154 ~| w4192;
assign w4242 = ~w4194;
assign w4243 = w4091 | w4195;
assign w4244 = w4172 | w4198;
assign w4245 = w4026 | w4201;
assign w4246 = w4111 ~^ w4202;
assign w4247 = w4168 ~^ w4203;
assign out1[4] = w4143 ~^ w4207;
assign w4248 = w4145 & w4207;
assign w4249 = w4190 ~^ w4208;
assign w4250 = w4190 | w4208;
assign w4251 = w4190 & w4208;
assign w4252 = w4183 | w4211;
assign w4253 = w4036 ~^ w4212;
assign w4254 = ~w4213;
assign w4255 = w4153 ~| w4215;
assign w4256 = w4095 ^ w4215;
assign w4257 = w4185 ~^ w4216;
assign w4258 = w4199 ~^ w4217;
assign w4259 = w4200 | w4217;
assign w4260 = w4196 ~^ w4218;
assign w4261 = ~w4218;
assign w4262 = w4219 & w4220;
assign w4263 = w3911 ~^ w4221;
assign w4264 = w3993 | w4222;
assign w4265 = w3648 | w4223;
assign w4266 = w4203 & w4224;
assign w4267 = w3974 ~| w4225;
assign w4268 = w4194 ~^ w4226;
assign w4269 = w4174 | w4228;
assign w4270 = w4182 & w4230;
assign w4271 = w4177 | w4231;
assign w4272 = w4180 | w4232;
assign w4273 = w4158 | w4236;
assign w4274 = w4024 | w4238;
assign w4275 = w4237 ~^ w4239;
assign w4276 = w4237 | w4239;
assign w4277 = w4237 & w4239;
assign w4278 = w4159 ~^ w4240;
assign w4279 = w4160 & w4240;
assign w4280 = w4193 | w4241;
assign w4281 = w4213 ~| w4242;
assign w4282 = w3974 ~^ w4247;
assign w4283 = w4144 | w4248;
assign w4284 = w4243 ~^ w4249;
assign w4285 = w4243 & w4250;
assign w4286 = w4214 & w4252;
assign w4287 = w4077 ~^ w4253;
assign w4288 = w4077 | w4253;
assign w4289 = w4077 & w4253;
assign w4290 = w4194 | w4254;
assign w4291 = w4152 | w4255;
assign w4292 = w4004 ~^ w4256;
assign w4293 = w4234 ~^ w4257;
assign w4294 = w4234 | w4257;
assign w4295 = w4234 & w4257;
assign w4296 = w4229 ~| w4258;
assign w4297 = w4229 & w4258;
assign w4298 = w4245 & w4259;
assign w4299 = ~w4260;
assign w4300 = w4197 | w4261;
assign w4301 = w4229 ^ w4262;
assign w4302 = w4264 & w4265;
assign w4303 = w4266 | w4267;
assign w4304 = w4213 ~^ w4268;
assign w4305 = w4209 ~^ w4269;
assign w4306 = w4149 & w4269;
assign w4307 = w4263 ~^ w4270;
assign w4308 = w4110 ~^ w4272;
assign w4309 = w4235 & w4273;
assign w4310 = w4161 | w4279;
assign w4311 = w4227 ~^ w4280;
assign w4312 = w4227 & w4280;
assign w4313 = w4227 | w4280;
assign w4314 = w4270 | w4282;
assign w4315 = w4270 & w4282;
assign out1[5] = w4204 ~^ w4283;
assign w4316 = w4206 & w4283;
assign w4317 = w4251 | w4285;
assign w4318 = w4226 & w4290;
assign w4319 = w4287 ~^ w4291;
assign w4320 = w4288 & w4291;
assign w4321 = w4284 & w4292;
assign w4322 = w4284 ~| w4292;
assign w4323 = w4286 ^ w4292;
assign w4324 = w4262 ~| w4297;
assign w4325 = w4189 ~| w4298;
assign w4326 = w4132 ^ w4298;
assign w4327 = w4244 & w4300;
assign w4328 = w4258 ~^ w4301;
assign w4329 = w3956 ^ w4302;
assign w4330 = w3956 ~| w4303;
assign w4331 = w3956 & w4303;
assign w4332 = w4274 ~^ w4305;
assign w4333 = ~w4305;
assign w4334 = w4210 | w4306;
assign w4335 = w4282 ~^ w4307;
assign w4336 = w4061 ~^ w4308;
assign w4337 = w4304 ~^ w4309;
assign w4338 = w4304 | w4309;
assign w4339 = w4304 & w4309;
assign w4340 = w4310 ~^ w4311;
assign w4341 = w4310 & w4313;
assign w4342 = w4263 | w4315;
assign w4343 = w4205 | w4316;
assign w4344 = w4281 | w4318;
assign w4345 = w4278 ~^ w4319;
assign w4346 = w4278 & w4319;
assign w4347 = w4278 | w4319;
assign w4348 = w4289 | w4320;
assign w4349 = w4286 ~| w4322;
assign w4350 = w4284 ~^ w4323;
assign w4351 = w4296 | w4324;
assign w4352 = w4188 | w4325;
assign w4353 = w4053 ~^ w4326;
assign w4354 = ~w4327;
assign w4355 = w4275 ~^ w4328;
assign w4356 = w4276 & w4328;
assign w4357 = w4303 ~^ w4329;
assign w4358 = w4302 ~| w4330;
assign w4359 = w4274 | w4333;
assign w4360 = w4274 & w4333;
assign w4361 = w4233 ~^ w4334;
assign w4362 = w4181 | w4334;
assign w4363 = ~w4334;
assign w4364 = w4271 ^ w4335;
assign w4365 = w4299 ~^ w4340;
assign w4366 = w4260 | w4340;
assign w4367 = ~w4340;
assign w4368 = w4312 | w4341;
assign w4369 = w4314 & w4342;
assign out1[6] = w4293 ~^ w4343;
assign w4370 = w4294 & w4343;
assign w4371 = ~w4344;
assign w4372 = w4317 ~^ w4345;
assign w4373 = w4317 & w4347;
assign w4374 = w4321 | w4349;
assign w4375 = w4344 ~^ w4350;
assign w4376 = w4344 ~| w4350;
assign w4377 = ~w4350;
assign w4378 = w4332 ~^ w4351;
assign w4379 = ~w4352;
assign w4380 = ~w4353;
assign w4381 = w4354 | w4355;
assign w4382 = ~w4355;
assign w4383 = w4277 | w4356;
assign w4384 = w4131 ~^ w4357;
assign w4385 = ~w4357;
assign w4386 = w4331 ~| w4358;
assign w4387 = w4351 & w4359;
assign w4388 = w4246 ~^ w4361;
assign w4389 = w4246 & w4362;
assign w4390 = w4233 ~| w4363;
assign w4391 = w4348 ~^ w4365;
assign w4392 = w4348 & w4366;
assign w4393 = w4299 ~| w4367;
assign w4394 = w4354 ~^ w4368;
assign w4395 = w4131 ~| w4369;
assign w4396 = w4131 & w4369;
assign w4397 = w4295 | w4370;
assign w4398 = ~w4372;
assign w4399 = w4346 | w4373;
assign w4400 = w4372 ~| w4374;
assign w4401 = ~w4374;
assign w4402 = w4371 | w4377;
assign w4403 = ~w4378;
assign w4404 = w4378 ~| w4380;
assign w4405 = w4368 & w4381;
assign w4406 = w4327 ~| w4382;
assign w4407 = w4369 ~^ w4384;
assign w4408 = w4336 ~^ w4386;
assign w4409 = w4360 | w4387;
assign w4410 = w4379 | w4388;
assign w4411 = ~w4388;
assign w4412 = w4389 | w4390;
assign w4413 = w4392 | w4393;
assign w4414 = w4382 ~^ w4394;
assign w4415 = w4385 ~| w4396;
assign out1[7] = w4337 ~^ w4397;
assign w4416 = ~w4397;
assign w4417 = w4374 ~^ w4398;
assign w4418 = w4391 ~^ w4399;
assign w4419 = ~w4399;
assign w4420 = w4398 | w4401;
assign w4421 = w4380 ~^ w4403;
assign w4422 = w4353 | w4403;
assign w4423 = w4405 | w4406;
assign w4424 = ~w4409;
assign w4425 = w4379 ~^ w4411;
assign w4426 = w4352 ~| w4411;
assign w4427 = w4364 ~^ w4412;
assign w4428 = w4271 ~| w4412;
assign w4429 = w4271 & w4412;
assign w4430 = ~w4413;
assign w4431 = ~w4414;
assign w4432 = w4395 ~| w4415;
assign w4433 = w4339 | w4416;
assign w4434 = w4391 & w4419;
assign w4435 = w4391 ~| w4419;
assign w4436 = w4383 ~^ w4421;
assign w4437 = w4383 & w4422;
assign w4438 = ~w4423;
assign w4439 = w4409 ~^ w4425;
assign w4440 = w4424 | w4426;
assign w4441 = ~w4427;
assign w4442 = w4335 ~| w4428;
assign w4443 = w4414 | w4430;
assign w4444 = w4413 ~^ w4431;
assign w4445 = w4413 ~| w4431;
assign w4446 = w4408 ~^ w4432;
assign w4447 = w4338 & w4433;
assign w4448 = w4423 ~^ w4436;
assign w4449 = w4404 | w4437;
assign w4450 = w4436 ~| w4438;
assign w4451 = w4436 & w4438;
assign w4452 = ~w4439;
assign w4453 = w4410 & w4440;
assign w4454 = w4429 | w4442;
assign w4455 = w4376 | w4447;
assign out1[8] = w4375 ^ w4447;
assign w4456 = ~w4449;
assign w4457 = w4449 ~^ w4452;
assign w4458 = w4449 ~| w4452;
assign w4459 = w4427 ~^ w4453;
assign w4460 = w4441 & w4453;
assign w4461 = w4441 ~| w4453;
assign w4462 = w4407 ~^ w4454;
assign w4463 = w4407 | w4454;
assign w4464 = w4407 & w4454;
assign w4465 = w4402 & w4455;
assign w4466 = w4439 | w4456;
assign out1[9] = w4417 ~^ w4465;
assign w4467 = w4400 | w4465;
assign w4468 = w4420 & w4467;
assign out1[10] = w4418 ~^ w4468;
assign w4469 = w4434 ~| w4468;
assign w4470 = w4435 | w4469;
assign out1[11] = w4444 ~^ w4470;
assign w4471 = ~w4470;
assign w4472 = w4445 | w4471;
assign w4473 = w4443 & w4472;
assign out1[12] = w4448 ~^ w4473;
assign w4474 = w4451 ~| w4473;
assign w4475 = w4450 | w4474;
assign out1[13] = w4457 ~^ w4475;
assign w4476 = ~w4475;
assign w4477 = w4458 | w4476;
assign w4478 = w4466 & w4477;
assign out1[14] = w4459 ~^ w4478;
assign w4479 = w4460 ~| w4478;
assign w4480 = w4461 | w4479;
assign out1[15] = w4462 ~^ w4480;
assign w4481 = w4463 & w4480;
assign w4482 = w4464 ~| w4481;
assign out1[16] = w4446 ~^ w4482;
wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482;
endmodule
module top(in1, in2, in3, out1, out2);
input wire [7:0] in1;
input wire [7:0] in2;
input wire [7:0] in3;
output wire [23:0] out1;
output wire [15:0] out2;

module top(in1, in2, in3, in4, out1, out2, out3, out4);
input wire [33:0] in1;
input wire [34:0] in2;
input wire [34:0] in3;
input wire [34:0] in4;
output wire out1;
output wire out2;
output wire out3;
output wire out4;
assign w0 = ~in1[0];
assign w1 = ~in1[0];
assign w2 = in1[1] & in1[0];
assign w3 = ~in1[1];
assign w4 = ~in1[2];
assign w5 = ~in1[3];
assign w6 = in1[5] ~| in1[4];
assign w7 = ~in1[6];
assign w8 = ~in1[7];
assign w9 = in1[9] | in1[8];
assign w10 = in1[13] ~| in1[12];
assign w11 = ~in1[14];
assign w12 = ~in1[15];
assign w13 = in1[17] | in1[16];
assign w14 = in1[21] | in1[20];
assign w15 = in1[23] | in1[22];
assign w16 = in1[25] | in1[24];
assign w17 = in1[29] ~| in1[28];
assign w18 = ~in1[30];
assign w19 = ~in1[31];
assign w20 = ~in1[32];
assign w21 = ~in1[33];
assign w22 = ~in2[0];
assign w23 = ~in2[1];
assign w24 = ~in2[4];
assign w25 = ~in2[22];
assign w26 = in1[0] ~^ in3[0];
assign w27 = in1[0] ~^ in4[0];
assign w28 = ~in4[2];
assign w29 = ~in4[16];
assign w30 = ~in4[18];
assign w31 = ~in4[21];
assign w32 = ~in4[28];
assign w33 = ~in4[30];
assign w34 = ~in4[31];
assign w35 = ~in4[33];
assign w36 = ~w0;
assign w37 = w1 & w3;
assign w38 = in1[11] | w9;
assign w39 = in1[19] | w13;
assign w40 = in1[27] | w16;
assign w41 = w0 | w22;
assign w42 = w36 | in4[0];
assign w43 = w4 & w37;
assign w44 = w2 | w37;
assign w45 = w37 ^ in1[2];
assign w46 = in1[10] ~| w38;
assign w47 = in1[18] | w39;
assign w48 = in1[26] ~| w40;
assign w49 = w23 | w41;
assign w50 = ~w41;
assign w51 = in4[1] & w42;
assign w52 = in4[1] ~| w42;
assign w53 = w5 & w43;
assign w54 = ~w43;
assign w55 = w44 ^ in4[1];
assign w56 = w44 ^ in3[1];
assign w57 = ~w45;
assign w58 = w45 ^ in4[2];
assign w59 = w45 ^ in3[2];
assign w60 = w28 ~| w45;
assign w61 = w28 & w45;
assign w62 = w14 | w47;
assign w63 = w44 & w49;
assign w64 = in2[1] ~| w50;
assign w65 = w44 ~| w52;
assign w66 = w6 & w53;
assign w67 = ~w53;
assign w68 = in1[3] & w54;
assign w69 = w27 | w55;
assign w70 = w26 | w56;
assign w71 = w57 ~| in2[2];
assign w72 = in2[2] & w57;
assign w73 = w15 ~| w62;
assign w74 = w63 ~| w64;
assign w75 = w51 ~| w65;
assign w76 = w7 & w66;
assign w77 = w66 ^ in1[6];
assign w78 = w67 ~^ in1[4];
assign w79 = in1[4] | w67;
assign w80 = w53 | w68;
assign w81 = w72 ~| w74;
assign w82 = w61 ~| w75;
assign w83 = w8 & w76;
assign w84 = ~w76;
assign w85 = ~w77;
assign w86 = ~w77;
assign w87 = w77 ^ in3[6];
assign w88 = w77 ^ in4[6];
assign w89 = ~w78;
assign w90 = w78 ^ in4[4];
assign w91 = w78 ^ in3[4];
assign w92 = w24 ~| w78;
assign w93 = w24 & w78;
assign w94 = w79 ~^ in1[5];
assign w95 = ~w80;
assign w96 = ~w80;
assign w97 = w80 ^ in4[3];
assign w98 = w80 ^ in3[3];
assign w99 = w71 ~| w81;
assign w100 = w60 ~| w82;
assign w101 = w46 & w83;
assign w102 = ~w83;
assign w103 = in1[7] & w84;
assign w104 = w85 ~| in4[6];
assign w105 = in4[6] & w85;
assign w106 = w86 ~| in2[6];
assign w107 = in2[6] & w86;
assign w108 = w89 ~| in4[4];
assign w109 = in4[4] & w89;
assign w110 = ~w94;
assign w111 = ~w94;
assign w112 = w94 ^ in3[5];
assign w113 = w94 ^ in4[5];
assign w114 = w95 ~| in4[3];
assign w115 = in4[3] & w95;
assign w116 = w96 ~| in2[3];
assign w117 = in2[3] & w96;
assign w118 = w58 | w97;
assign w119 = w59 | w98;
assign w120 = w10 & w101;
assign w121 = ~w101;
assign w122 = w102 ~^ in1[8];
assign w123 = in1[8] | w102;
assign w124 = w9 | w102;
assign w125 = w83 | w103;
assign w126 = w110 ~| in4[5];
assign w127 = in4[5] & w110;
assign w128 = w111 ~| in2[5];
assign w129 = in2[5] & w111;
assign w130 = w91 | w112;
assign w131 = w90 | w113;
assign w132 = w100 ~| w114;
assign w133 = w99 ~| w117;
assign w134 = w69 | w118;
assign w135 = w70 | w119;
assign w136 = w11 & w120;
assign w137 = w120 ^ in1[14];
assign w138 = w121 ~^ in1[12];
assign w139 = in1[12] | w121;
assign w140 = ~w122;
assign w141 = ~w122;
assign w142 = w122 ^ in4[8];
assign w143 = w122 ^ in3[8];
assign w144 = w123 ~^ in1[9];
assign w145 = w124 ~^ in1[10];
assign w146 = in1[10] | w124;
assign w147 = ~w125;
assign w148 = ~w125;
assign w149 = w125 ^ in3[7];
assign w150 = w125 ^ in4[7];
assign w151 = w115 ~| w132;
assign w152 = w116 ~| w133;
assign w153 = w12 & w136;
assign w154 = w12 ~| w136;
assign w155 = ~w137;
assign w156 = ~w137;
assign w157 = w137 ^ in4[14];
assign w158 = w137 ^ in3[14];
assign w159 = ~w138;
assign w160 = ~w138;
assign w161 = w138 ^ in3[12];
assign w162 = w138 ^ in4[12];
assign w163 = w139 ~^ in1[13];
assign w164 = w140 ~| in4[8];
assign w165 = in4[8] & w140;
assign w166 = w141 ~| in2[8];
assign w167 = in2[8] & w141;
assign w168 = ~w144;
assign w169 = ~w144;
assign w170 = w144 ^ in3[9];
assign w171 = w144 ^ in4[9];
assign w172 = ~w145;
assign w173 = ~w145;
assign w174 = w145 ^ in3[10];
assign w175 = w145 ^ in4[10];
assign w176 = w146 ~^ in1[11];
assign w177 = w147 ~| in4[7];
assign w178 = in4[7] & w147;
assign w179 = w148 ~| in2[7];
assign w180 = in2[7] & w148;
assign w181 = w87 | w149;
assign w182 = w88 | w150;
assign w183 = w108 ~| w151;
assign w184 = w92 ~| w152;
assign w185 = w73 & w153;
assign w186 = ~w153;
assign w187 = ~w153;
assign w188 = w153 | w154;
assign w189 = w155 ~| in4[14];
assign w190 = in4[14] & w155;
assign w191 = w156 ~| in2[14];
assign w192 = in2[14] & w156;
assign w193 = w159 ~| in4[12];
assign w194 = in4[12] & w159;
assign w195 = w160 ~| in2[12];
assign w196 = in2[12] & w160;
assign w197 = ~w163;
assign w198 = ~w163;
assign w199 = w163 ^ in3[13];
assign w200 = w163 ^ in4[13];
assign w201 = w168 ~| in4[9];
assign w202 = in4[9] & w168;
assign w203 = w169 ~| in2[9];
assign w204 = in2[9] & w169;
assign w205 = w143 | w170;
assign w206 = w142 | w171;
assign w207 = w172 ~| in4[10];
assign w208 = in4[10] & w172;
assign w209 = w173 ~| in2[10];
assign w210 = in2[10] & w173;
assign w211 = ~w176;
assign w212 = ~w176;
assign w213 = w176 ^ in3[11];
assign w214 = w176 ^ in4[11];
assign w215 = w130 | w181;
assign w216 = w131 | w182;
assign w217 = w109 ~| w183;
assign w218 = w93 ~| w184;
assign w219 = w48 & w185;
assign w220 = ~w185;
assign w221 = w185 ^ in1[24];
assign w222 = in1[16] | w186;
assign w223 = w13 | w186;
assign w224 = w187 ~^ in1[16];
assign w225 = w47 | w187;
assign w226 = ~w188;
assign w227 = ~w188;
assign w228 = w188 ^ in4[15];
assign w229 = w188 ^ in3[15];
assign w230 = w197 ~| in4[13];
assign w231 = in4[13] & w197;
assign w232 = w198 ~| in2[13];
assign w233 = in2[13] & w198;
assign w234 = w161 | w199;
assign w235 = w162 | w200;
assign w236 = w211 ~| in4[11];
assign w237 = in4[11] & w211;
assign w238 = w212 ~| in2[11];
assign w239 = in2[11] & w212;
assign w240 = w174 | w213;
assign w241 = w175 | w214;
assign w242 = w135 | w215;
assign w243 = w134 | w216;
assign w244 = w126 ~| w217;
assign w245 = w129 ~| w218;
assign w246 = w17 & w219;
assign w247 = ~w219;
assign w248 = w16 | w220;
assign w249 = in1[24] | w220;
assign w250 = ~w221;
assign w251 = ~w221;
assign w252 = w221 ^ in3[24];
assign w253 = w221 ^ in4[24];
assign w254 = w222 ~^ in1[17];
assign w255 = w223 ~^ in1[18];
assign w256 = in1[18] | w223;
assign w257 = ~w224;
assign w258 = w224 ^ in4[16];
assign w259 = w224 ^ in3[16];
assign w260 = w29 ~| w224;
assign w261 = w29 & w224;
assign w262 = w225 ~^ in1[20];
assign w263 = w14 | w225;
assign w264 = in1[20] | w225;
assign w265 = w226 ~| in4[15];
assign w266 = in4[15] & w226;
assign w267 = w227 ~| in2[15];
assign w268 = in2[15] & w227;
assign w269 = w157 | w228;
assign w270 = w158 | w229;
assign w271 = w205 | w240;
assign w272 = w206 | w241;
assign w273 = w127 ~| w244;
assign w274 = w128 ~| w245;
assign w275 = w18 & w246;
assign w276 = ~w246;
assign w277 = w247 ~^ in1[28];
assign w278 = in1[28] | w247;
assign w279 = w248 ~^ in1[26];
assign w280 = in1[26] | w248;
assign w281 = w249 ~^ in1[25];
assign w282 = w250 ~| in4[24];
assign w283 = in4[24] & w250;
assign w284 = w251 ~| in2[24];
assign w285 = in2[24] & w251;
assign w286 = ~w254;
assign w287 = ~w254;
assign w288 = w254 ^ in4[17];
assign w289 = w254 ^ in3[17];
assign w290 = ~w255;
assign w291 = w255 ^ in4[18];
assign w292 = w255 ^ in3[18];
assign w293 = w30 ~| w255;
assign w294 = w30 & w255;
assign w295 = w256 ~^ in1[19];
assign w296 = w257 ~| in2[16];
assign w297 = in2[16] & w257;
assign w298 = ~w262;
assign w299 = ~w262;
assign w300 = w262 ^ in4[20];
assign w301 = w262 ^ in3[20];
assign w302 = w263 ~^ in1[22];
assign w303 = in1[22] | w263;
assign w304 = w264 ~^ in1[21];
assign w305 = w235 | w269;
assign w306 = w234 | w270;
assign w307 = w104 ~| w273;
assign w308 = w107 ~| w274;
assign w309 = w19 & w275;
assign w310 = w275 ^ in1[31];
assign w311 = in1[30] & w276;
assign w312 = ~w277;
assign w313 = w277 ^ in4[28];
assign w314 = w277 ^ in3[28];
assign w315 = w32 ~| w277;
assign w316 = w32 & w277;
assign w317 = w278 ~^ in1[29];
assign w318 = ~w279;
assign w319 = ~w279;
assign w320 = w279 ^ in3[26];
assign w321 = w279 ^ in4[26];
assign w322 = w280 ~^ in1[27];
assign w323 = ~w281;
assign w324 = ~w281;
assign w325 = w281 ^ in3[25];
assign w326 = w281 ^ in4[25];
assign w327 = w286 ~| in4[17];
assign w328 = in4[17] & w286;
assign w329 = w287 ~| in2[17];
assign w330 = in2[17] & w287;
assign w331 = w258 | w288;
assign w332 = w259 | w289;
assign w333 = w290 ~| in2[18];
assign w334 = in2[18] & w290;
assign w335 = ~w295;
assign w336 = ~w295;
assign w337 = w295 ^ in4[19];
assign w338 = w295 ^ in3[19];
assign w339 = w298 ~| in4[20];
assign w340 = in4[20] & w298;
assign w341 = w299 ~| in2[20];
assign w342 = in2[20] & w299;
assign w343 = ~w302;
assign w344 = w302 ^ in4[22];
assign w345 = w302 ^ in3[22];
assign w346 = w25 ~| w302;
assign w347 = w25 & w302;
assign w348 = w303 ~^ in1[23];
assign w349 = ~w304;
assign w350 = w304 ^ in3[21];
assign w351 = w304 ^ in4[21];
assign w352 = w31 ~| w304;
assign w353 = w31 & w304;
assign w354 = w272 | w305;
assign w355 = w271 | w306;
assign w356 = w105 ~| w307;
assign w357 = w106 ~| w308;
assign w358 = w20 & w309;
assign w359 = ~w309;
assign w360 = ~w310;
assign w361 = w310 ^ in3[31];
assign w362 = w310 ^ in4[31];
assign w363 = w34 ~| w310;
assign w364 = w34 & w310;
assign w365 = w275 | w311;
assign w366 = w312 ~| in2[28];
assign w367 = in2[28] & w312;
assign w368 = ~w317;
assign w369 = ~w317;
assign w370 = w317 ^ in3[29];
assign w371 = w317 ^ in4[29];
assign w372 = w318 ~| in4[26];
assign w373 = in4[26] & w318;
assign w374 = w319 ~| in2[26];
assign w375 = in2[26] & w319;
assign w376 = ~w322;
assign w377 = ~w322;
assign w378 = w322 ^ in3[27];
assign w379 = w322 ^ in4[27];
assign w380 = w323 ~| in4[25];
assign w381 = in4[25] & w323;
assign w382 = w324 ~| in2[25];
assign w383 = in2[25] & w324;
assign w384 = w252 | w325;
assign w385 = w253 | w326;
assign w386 = w335 ~| in4[19];
assign w387 = in4[19] & w335;
assign w388 = w336 ~| in2[19];
assign w389 = in2[19] & w336;
assign w390 = w291 | w337;
assign w391 = w292 | w338;
assign w392 = w343 ~| in4[22];
assign w393 = in4[22] & w343;
assign w394 = ~w348;
assign w395 = ~w348;
assign w396 = w348 ^ in3[23];
assign w397 = w348 ^ in4[23];
assign w398 = w349 ~| in2[21];
assign w399 = in2[21] & w349;
assign w400 = w301 | w350;
assign w401 = w300 | w351;
assign w402 = w243 | w354;
assign w403 = w242 | w355;
assign w404 = w177 ~| w356;
assign w405 = w180 ~| w357;
assign w406 = w21 & w358;
assign w407 = w358 ^ in1[33];
assign w408 = in1[32] & w359;
assign w409 = w360 ~| in2[31];
assign w410 = in2[31] & w360;
assign w411 = ~w365;
assign w412 = w365 ^ in3[30];
assign w413 = w365 ^ in4[30];
assign w414 = w33 ~| w365;
assign w415 = w33 & w365;
assign w416 = w368 ~| in4[29];
assign w417 = in4[29] & w368;
assign w418 = w369 ~| in2[29];
assign w419 = in2[29] & w369;
assign w420 = w314 | w370;
assign w421 = w313 | w371;
assign w422 = w376 ~| in4[27];
assign w423 = in4[27] & w376;
assign w424 = w377 ~| in2[27];
assign w425 = in2[27] & w377;
assign w426 = w320 | w378;
assign w427 = w321 | w379;
assign w428 = w331 | w390;
assign w429 = w332 | w391;
assign w430 = w394 ~| in4[23];
assign w431 = in4[23] & w394;
assign w432 = w395 ~| in2[23];
assign w433 = in2[23] & w395;
assign w434 = w345 | w396;
assign w435 = w344 | w397;
assign w436 = w178 ~| w404;
assign w437 = w179 ~| w405;
assign w438 = ~w407;
assign w439 = w407 ^ in4[33];
assign w440 = w407 ^ in3[33];
assign w441 = w35 ~| w407;
assign w442 = w35 & w407;
assign w443 = w358 | w408;
assign w444 = w411 ~| in2[30];
assign w445 = in2[30] & w411;
assign w446 = w361 | w412;
assign w447 = w362 | w413;
assign w448 = w384 | w426;
assign w449 = w385 | w427;
assign w450 = w400 | w434;
assign w451 = w401 | w435;
assign w452 = w164 ~| w436;
assign w453 = w167 ~| w437;
assign w454 = w438 ~| in2[33];
assign w455 = in2[33] & w438;
assign w456 = ~w443;
assign w457 = ~w443;
assign w458 = w443 ^ in4[32];
assign w459 = w443 ^ in3[32];
assign w460 = w420 | w446;
assign w461 = w421 | w447;
assign w462 = w429 | w450;
assign w463 = w428 | w451;
assign w464 = w165 ~| w452;
assign w465 = w166 ~| w453;
assign w466 = w456 ~| in4[32];
assign w467 = in4[32] & w456;
assign w468 = w457 ~| in2[32];
assign w469 = in2[32] & w457;
assign w470 = w439 | w458;
assign w471 = w448 | w460;
assign w472 = w449 | w461;
assign w473 = w201 ~| w464;
assign w474 = w204 ~| w465;
assign w475 = w202 ~| w473;
assign w476 = w203 ~| w474;
assign w477 = w207 ~| w475;
assign w478 = w210 ~| w476;
assign w479 = w208 ~| w477;
assign w480 = w209 ~| w478;
assign w481 = w236 ~| w479;
assign w482 = w239 ~| w480;
assign w483 = w237 ~| w481;
assign w484 = w238 ~| w482;
assign w485 = w193 ~| w483;
assign w486 = w196 ~| w484;
assign w487 = w194 ~| w485;
assign w488 = w195 ~| w486;
assign w489 = w230 ~| w487;
assign w490 = w233 ~| w488;
assign w491 = w231 ~| w489;
assign w492 = w232 ~| w490;
assign w493 = w189 ~| w491;
assign w494 = w192 ~| w492;
assign w495 = w190 ~| w493;
assign w496 = w191 ~| w494;
assign w497 = w265 ~| w495;
assign w498 = w268 ~| w496;
assign w499 = w266 ~| w497;
assign w500 = w267 ~| w498;
assign w501 = w261 ~| w499;
assign w502 = w297 ~| w500;
assign w503 = w260 ~| w501;
assign w504 = w296 ~| w502;
assign w505 = w327 ~| w503;
assign w506 = w330 ~| w504;
assign w507 = w328 ~| w505;
assign w508 = w329 ~| w506;
assign w509 = w294 ~| w507;
assign w510 = w334 ~| w508;
assign w511 = w293 ~| w509;
assign w512 = w333 ~| w510;
assign w513 = w386 ~| w511;
assign w514 = w389 ~| w512;
assign w515 = w387 ~| w513;
assign w516 = w388 ~| w514;
assign w517 = w339 ~| w515;
assign w518 = w342 ~| w516;
assign w519 = w340 ~| w517;
assign w520 = w341 ~| w518;
assign w521 = w353 ~| w519;
assign w522 = w399 ~| w520;
assign w523 = w352 ~| w521;
assign w524 = w398 ~| w522;
assign w525 = w392 ~| w523;
assign w526 = w346 ~| w524;
assign w527 = w393 ~| w525;
assign w528 = w347 ~| w526;
assign w529 = w430 ~| w527;
assign w530 = w433 ~| w528;
assign w531 = w431 ~| w529;
assign w532 = w432 ~| w530;
assign w533 = w282 ~| w531;
assign w534 = w285 ~| w532;
assign w535 = w283 ~| w533;
assign w536 = w284 ~| w534;
assign w537 = w380 ~| w535;
assign w538 = w383 ~| w536;
assign w539 = w381 ~| w537;
assign w540 = w382 ~| w538;
assign w541 = w372 ~| w539;
assign w542 = w375 ~| w540;
assign w543 = w373 ~| w541;
assign w544 = w374 ~| w542;
assign w545 = w422 ~| w543;
assign w546 = w425 ~| w544;
assign w547 = w423 ~| w545;
assign w548 = w424 ~| w546;
assign w549 = w316 ~| w547;
assign w550 = w367 ~| w548;
assign w551 = w315 ~| w549;
assign w552 = w366 ~| w550;
assign w553 = w416 ~| w551;
assign w554 = w419 ~| w552;
assign w555 = w417 ~| w553;
assign w556 = w418 ~| w554;
assign w557 = w415 ~| w555;
assign w558 = w445 ~| w556;
assign w559 = w414 ~| w557;
assign w560 = w444 ~| w558;
assign w561 = w364 ~| w559;
assign w562 = w410 ~| w560;
assign w563 = w363 ~| w561;
assign w564 = w409 ~| w562;
assign w565 = w466 ~| w563;
assign w566 = w469 ~| w564;
assign w567 = w467 ~| w565;
assign w568 = w468 ~| w566;
assign w569 = w442 ~| w567;
assign w570 = w455 ~| w568;
assign w571 = w441 | w569;
assign w572 = w454 ~| w570;
assign w573 = w406 ~| w572;
assign out1 = in2[34] | w573;
wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573;
endmodule
module top(in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, out1);
input wire [8:0] in1;
input wire in10;
input wire in11;
input wire [8:0] in12;
input wire [7:0] in13;
input wire in14;
input wire in15;
input wire [8:0] in16;
input wire [7:0] in17;
input wire in18;
input wire in19;
input wire [7:0] in2;
input wire [8:0] in20;
input wire [7:0] in21;
input wire in22;
input wire in23;
input wire [8:0] in24;
input wire [7:0] in25;
input wire in3;
input wire in4;
input wire [6:0] in5;
input wire in6;
input wire in7;
input wire [8:0] in8;
input wire [7:0] in9;
output wire [16:0] out1;
assign w0 = ~in10;
assign w1 = ~in10;
assign w2 = ~in10;
assign w3 = ~in10;
assign w4 = ~in10;
assign w5 = ~in10;
assign w6 = ~in10;
assign w7 = ~in10;
assign w8 = ~in10;
assign w9 = ~in10;
assign w10 = ~in10;
assign w11 = ~in10;
assign w12 = ~in10;
assign w13 = ~in10;
assign w14 = ~in10;
assign w15 = ~in10;
assign w16 = ~in12[0];
assign w17 = ~in12[0];
assign w18 = ~in12[0];
assign w19 = ~in12[0];
assign w20 = ~in12[1];
assign w21 = ~in12[1];
assign w22 = ~in12[1];
assign w23 = ~in12[1];
assign w24 = ~in12[2];
assign w25 = ~in12[3];
assign w26 = ~in12[4];
assign w27 = ~in12[5];
assign w28 = ~in12[6];
assign w29 = ~in12[7];
assign w30 = ~in12[8];
assign w31 = in12[5] & in13[0];
assign w32 = in12[3] & in13[0];
assign w33 = in12[4] & in13[0];
assign w34 = in12[6] & in13[0];
assign w35 = ~in13[0];
assign w36 = in12[8] & in13[1];
assign w37 = in12[4] & in13[1];
assign w38 = ~in13[1];
assign w39 = ~in13[1];
assign w40 = ~in13[1];
assign w41 = ~in13[1];
assign w42 = in12[7] & in13[2];
assign w43 = ~in13[2];
assign w44 = ~in13[2];
assign w45 = ~in13[2];
assign w46 = ~in13[2];
assign w47 = ~in13[3];
assign w48 = ~in13[3];
assign w49 = ~in13[3];
assign w50 = ~in13[3];
assign w51 = ~in13[3];
assign w52 = ~in13[4];
assign w53 = ~in13[4];
assign w54 = ~in13[4];
assign w55 = ~in13[4];
assign w56 = ~in13[4];
assign w57 = in12[3] & in13[5];
assign w58 = in12[0] & in13[5];
assign w59 = ~in13[5];
assign w60 = in12[2] & in13[6];
assign w61 = ~in13[6];
assign w62 = ~in13[6];
assign w63 = ~in13[6];
assign w64 = ~in13[6];
assign w65 = in12[8] & in13[7];
assign w66 = ~in13[7];
assign w67 = ~in13[7];
assign w68 = ~in13[7];
assign w69 = ~in13[7];
assign w70 = ~in14;
assign w71 = ~in14;
assign w72 = ~in14;
assign w73 = ~in14;
assign w74 = ~in14;
assign w75 = ~in14;
assign w76 = ~in14;
assign w77 = ~in14;
assign w78 = ~in14;
assign w79 = ~in14;
assign w80 = ~in14;
assign w81 = ~in14;
assign w82 = ~in14;
assign w83 = ~in14;
assign w84 = ~in14;
assign w85 = ~in14;
assign w86 = ~in16[0];
assign w87 = ~in16[0];
assign w88 = ~in16[0];
assign w89 = ~in16[0];
assign w90 = ~in16[1];
assign w91 = ~in16[1];
assign w92 = ~in16[1];
assign w93 = ~in16[1];
assign w94 = ~in16[2];
assign w95 = ~in16[3];
assign w96 = ~in16[4];
assign w97 = ~in16[5];
assign w98 = ~in16[6];
assign w99 = ~in16[7];
assign w100 = ~in16[8];
assign w101 = in16[5] & in17[0];
assign w102 = in16[3] & in17[0];
assign w103 = in16[4] & in17[0];
assign w104 = in16[6] & in17[0];
assign w105 = ~in17[0];
assign w106 = in16[8] & in17[1];
assign w107 = in16[4] & in17[1];
assign w108 = ~in17[1];
assign w109 = ~in17[1];
assign w110 = ~in17[1];
assign w111 = ~in17[1];
assign w112 = in16[7] & in17[2];
assign w113 = ~in17[2];
assign w114 = ~in17[2];
assign w115 = ~in17[2];
assign w116 = ~in17[2];
assign w117 = ~in17[3];
assign w118 = ~in17[3];
assign w119 = ~in17[3];
assign w120 = ~in17[3];
assign w121 = ~in17[3];
assign w122 = ~in17[4];
assign w123 = ~in17[4];
assign w124 = ~in17[4];
assign w125 = ~in17[4];
assign w126 = ~in17[4];
assign w127 = in16[3] & in17[5];
assign w128 = in16[0] & in17[5];
assign w129 = ~in17[5];
assign w130 = in16[2] & in17[6];
assign w131 = ~in17[6];
assign w132 = ~in17[6];
assign w133 = ~in17[6];
assign w134 = ~in17[6];
assign w135 = in16[8] & in17[7];
assign w136 = ~in17[7];
assign w137 = ~in17[7];
assign w138 = ~in17[7];
assign w139 = ~in17[7];
assign w140 = ~in18;
assign w141 = ~in18;
assign w142 = ~in18;
assign w143 = ~in18;
assign w144 = ~in18;
assign w145 = ~in18;
assign w146 = ~in18;
assign w147 = ~in18;
assign w148 = ~in18;
assign w149 = ~in18;
assign w150 = ~in18;
assign w151 = ~in18;
assign w152 = ~in18;
assign w153 = ~in18;
assign w154 = ~in18;
assign w155 = ~in18;
assign w156 = ~in1[0];
assign w157 = ~in1[0];
assign w158 = ~in1[0];
assign w159 = ~in1[0];
assign w160 = ~in1[1];
assign w161 = ~in1[1];
assign w162 = ~in1[1];
assign w163 = ~in1[1];
assign w164 = ~in1[2];
assign w165 = ~in1[3];
assign w166 = ~in1[4];
assign w167 = ~in1[5];
assign w168 = ~in1[6];
assign w169 = ~in1[7];
assign w170 = ~in1[8];
assign w171 = ~in20[0];
assign w172 = ~in20[0];
assign w173 = ~in20[0];
assign w174 = ~in20[0];
assign w175 = ~in20[1];
assign w176 = ~in20[1];
assign w177 = ~in20[1];
assign w178 = ~in20[1];
assign w179 = ~in20[2];
assign w180 = ~in20[3];
assign w181 = ~in20[4];
assign w182 = ~in20[5];
assign w183 = ~in20[6];
assign w184 = ~in20[7];
assign w185 = ~in20[8];
assign w186 = in20[5] & in21[0];
assign w187 = in20[3] & in21[0];
assign w188 = in20[4] & in21[0];
assign w189 = in20[6] & in21[0];
assign w190 = ~in21[0];
assign w191 = in20[8] & in21[1];
assign w192 = in20[4] & in21[1];
assign w193 = ~in21[1];
assign w194 = ~in21[1];
assign w195 = ~in21[1];
assign w196 = ~in21[1];
assign w197 = in20[7] & in21[2];
assign w198 = ~in21[2];
assign w199 = ~in21[2];
assign w200 = ~in21[2];
assign w201 = ~in21[2];
assign w202 = ~in21[3];
assign w203 = ~in21[3];
assign w204 = ~in21[3];
assign w205 = ~in21[3];
assign w206 = ~in21[3];
assign w207 = ~in21[4];
assign w208 = ~in21[4];
assign w209 = ~in21[4];
assign w210 = ~in21[4];
assign w211 = ~in21[4];
assign w212 = in20[3] & in21[5];
assign w213 = in20[0] & in21[5];
assign w214 = ~in21[5];
assign w215 = in20[2] & in21[6];
assign w216 = ~in21[6];
assign w217 = ~in21[6];
assign w218 = ~in21[6];
assign w219 = ~in21[6];
assign w220 = in20[8] & in21[7];
assign w221 = ~in21[7];
assign w222 = ~in21[7];
assign w223 = ~in21[7];
assign w224 = ~in21[7];
assign w225 = ~in22;
assign w226 = ~in22;
assign w227 = ~in22;
assign w228 = ~in22;
assign w229 = ~in22;
assign w230 = ~in22;
assign w231 = ~in22;
assign w232 = ~in22;
assign w233 = ~in22;
assign w234 = ~in22;
assign w235 = ~in22;
assign w236 = ~in22;
assign w237 = ~in22;
assign w238 = ~in22;
assign w239 = ~in22;
assign w240 = ~in22;
assign w241 = ~in24[0];
assign w242 = ~in24[0];
assign w243 = ~in24[0];
assign w244 = ~in24[0];
assign w245 = ~in24[1];
assign w246 = ~in24[1];
assign w247 = ~in24[1];
assign w248 = ~in24[1];
assign w249 = ~in24[2];
assign w250 = ~in24[3];
assign w251 = ~in24[4];
assign w252 = ~in24[5];
assign w253 = ~in24[6];
assign w254 = ~in24[7];
assign w255 = ~in24[8];
assign w256 = in24[5] & in25[0];
assign w257 = in24[3] & in25[0];
assign w258 = in24[4] & in25[0];
assign w259 = in24[6] & in25[0];
assign w260 = ~in25[0];
assign w261 = in24[8] & in25[1];
assign w262 = in24[4] & in25[1];
assign w263 = ~in25[1];
assign w264 = ~in25[1];
assign w265 = ~in25[1];
assign w266 = ~in25[1];
assign w267 = in24[7] & in25[2];
assign w268 = ~in25[2];
assign w269 = ~in25[2];
assign w270 = ~in25[2];
assign w271 = ~in25[2];
assign w272 = ~in25[3];
assign w273 = ~in25[3];
assign w274 = ~in25[3];
assign w275 = ~in25[3];
assign w276 = ~in25[3];
assign w277 = ~in25[4];
assign w278 = ~in25[4];
assign w279 = ~in25[4];
assign w280 = ~in25[4];
assign w281 = ~in25[4];
assign w282 = in24[3] & in25[5];
assign w283 = in24[0] & in25[5];
assign w284 = ~in25[5];
assign w285 = in24[2] & in25[6];
assign w286 = ~in25[6];
assign w287 = ~in25[6];
assign w288 = ~in25[6];
assign w289 = ~in25[6];
assign w290 = in24[8] & in25[7];
assign w291 = ~in25[7];
assign w292 = ~in25[7];
assign w293 = ~in25[7];
assign w294 = ~in25[7];
assign w295 = in1[5] & in2[0];
assign w296 = in1[3] & in2[0];
assign w297 = in1[4] & in2[0];
assign w298 = in1[6] & in2[0];
assign w299 = ~in2[0];
assign w300 = in1[8] & in2[1];
assign w301 = in1[4] & in2[1];
assign w302 = ~in2[1];
assign w303 = ~in2[1];
assign w304 = ~in2[1];
assign w305 = ~in2[1];
assign w306 = in1[7] & in2[2];
assign w307 = ~in2[2];
assign w308 = ~in2[2];
assign w309 = ~in2[2];
assign w310 = ~in2[2];
assign w311 = ~in2[3];
assign w312 = ~in2[3];
assign w313 = ~in2[3];
assign w314 = ~in2[3];
assign w315 = ~in2[3];
assign w316 = ~in2[4];
assign w317 = ~in2[4];
assign w318 = ~in2[4];
assign w319 = ~in2[4];
assign w320 = ~in2[4];
assign w321 = in1[3] & in2[5];
assign w322 = in1[0] & in2[5];
assign w323 = ~in2[5];
assign w324 = in1[2] & in2[6];
assign w325 = ~in2[6];
assign w326 = ~in2[6];
assign w327 = ~in2[6];
assign w328 = ~in2[6];
assign w329 = in1[8] & in2[7];
assign w330 = ~in2[7];
assign w331 = ~in2[7];
assign w332 = ~in2[7];
assign w333 = ~in2[7];
assign w334 = ~in3;
assign w335 = ~in3;
assign w336 = ~in3;
assign w337 = ~in3;
assign w338 = ~in3;
assign w339 = ~in3;
assign w340 = ~in3;
assign w341 = ~in3;
assign w342 = ~in3;
assign w343 = ~in3;
assign w344 = ~in3;
assign w345 = ~in3;
assign w346 = ~in3;
assign w347 = ~in3;
assign w348 = ~in3;
assign w349 = ~in3;
assign w350 = ~in5[1];
assign w351 = ~in5[2];
assign w352 = ~in5[3];
assign w353 = ~in6;
assign w354 = ~in6;
assign w355 = ~in6;
assign w356 = ~in6;
assign w357 = ~in6;
assign w358 = ~in6;
assign w359 = ~in6;
assign w360 = ~in6;
assign w361 = ~in6;
assign w362 = ~in6;
assign w363 = ~in6;
assign w364 = ~in6;
assign w365 = ~in6;
assign w366 = ~in6;
assign w367 = ~in6;
assign w368 = ~in6;
assign w369 = ~in8[0];
assign w370 = ~in8[0];
assign w371 = ~in8[0];
assign w372 = ~in8[0];
assign w373 = ~in8[1];
assign w374 = ~in8[1];
assign w375 = ~in8[1];
assign w376 = ~in8[1];
assign w377 = ~in8[2];
assign w378 = ~in8[3];
assign w379 = ~in8[4];
assign w380 = ~in8[5];
assign w381 = ~in8[6];
assign w382 = ~in8[7];
assign w383 = ~in8[8];
assign w384 = in8[5] & in9[0];
assign w385 = in8[3] & in9[0];
assign w386 = in8[4] & in9[0];
assign w387 = in8[6] & in9[0];
assign w388 = ~in9[0];
assign w389 = in8[8] & in9[1];
assign w390 = in8[4] & in9[1];
assign w391 = ~in9[1];
assign w392 = ~in9[1];
assign w393 = ~in9[1];
assign w394 = ~in9[1];
assign w395 = in8[7] & in9[2];
assign w396 = ~in9[2];
assign w397 = ~in9[2];
assign w398 = ~in9[2];
assign w399 = ~in9[2];
assign w400 = ~in9[3];
assign w401 = ~in9[3];
assign w402 = ~in9[3];
assign w403 = ~in9[3];
assign w404 = ~in9[3];
assign w405 = ~in9[4];
assign w406 = ~in9[4];
assign w407 = ~in9[4];
assign w408 = ~in9[4];
assign w409 = ~in9[4];
assign w410 = in8[3] & in9[5];
assign w411 = in8[0] & in9[5];
assign w412 = ~in9[5];
assign w413 = in8[2] & in9[6];
assign w414 = ~in9[6];
assign w415 = ~in9[6];
assign w416 = ~in9[6];
assign w417 = ~in9[6];
assign w418 = in8[8] & in9[7];
assign w419 = ~in9[7];
assign w420 = ~in9[7];
assign w421 = ~in9[7];
assign w422 = ~in9[7];
assign w423 = w24 | w35;
assign w424 = w18 ~| w35;
assign w425 = w20 ~| w35;
assign w426 = w30 | w35;
assign w427 = w29 | w35;
assign w428 = w31 & w37;
assign w429 = w31 ~^ w37;
assign w430 = w16 ~| w38;
assign w431 = w29 | w38;
assign w432 = w28 | w39;
assign w433 = w25 | w39;
assign w434 = w22 ~| w40;
assign w435 = w24 | w41;
assign w436 = w27 | w41;
assign w437 = w36 & w42;
assign w438 = w36 ~^ w42;
assign w439 = w26 | w43;
assign w440 = w25 | w43;
assign w441 = w27 | w44;
assign w442 = w19 | w44;
assign w443 = w24 | w45;
assign w444 = w30 | w45;
assign w445 = w28 | w46;
assign w446 = w20 | w46;
assign w447 = w27 | w47;
assign w448 = w30 | w47;
assign w449 = w24 | w48;
assign w450 = w26 | w48;
assign w451 = w28 | w49;
assign w452 = w17 | w49;
assign w453 = w22 | w50;
assign w454 = w29 | w50;
assign w455 = w25 | w51;
assign w456 = w26 | w52;
assign w457 = w30 | w52;
assign w458 = w27 | w53;
assign w459 = w29 | w53;
assign w460 = w24 | w54;
assign w461 = w28 | w54;
assign w462 = w21 | w55;
assign w463 = w25 | w55;
assign w464 = w19 | w56;
assign w465 = ~w57;
assign w466 = ~w58;
assign w467 = w27 | w59;
assign w468 = w23 | w59;
assign w469 = w30 | w59;
assign w470 = w26 | w59;
assign w471 = w24 | w59;
assign w472 = w29 | w59;
assign w473 = w28 | w59;
assign w474 = w57 | w60;
assign w475 = ~w60;
assign w476 = w27 | w61;
assign w477 = w29 | w61;
assign w478 = w26 | w62;
assign w479 = w17 | w62;
assign w480 = w25 | w63;
assign w481 = w23 | w63;
assign w482 = w30 | w64;
assign w483 = w28 | w64;
assign w484 = w5 & w65;
assign w485 = w27 | w66;
assign w486 = w26 | w66;
assign w487 = w29 | w67;
assign w488 = w21 | w67;
assign w489 = w28 | w68;
assign w490 = w24 | w68;
assign w491 = w25 | w69;
assign w492 = w16 | w69;
assign w493 = w94 | w105;
assign w494 = w88 ~| w105;
assign w495 = w90 ~| w105;
assign w496 = w100 | w105;
assign w497 = w99 | w105;
assign w498 = w101 & w107;
assign w499 = w101 ~^ w107;
assign w500 = w86 ~| w108;
assign w501 = w99 | w108;
assign w502 = w98 | w109;
assign w503 = w95 | w109;
assign w504 = w92 ~| w110;
assign w505 = w94 | w111;
assign w506 = w97 | w111;
assign w507 = w106 & w112;
assign w508 = w106 ~^ w112;
assign w509 = w96 | w113;
assign w510 = w95 | w113;
assign w511 = w97 | w114;
assign w512 = w89 | w114;
assign w513 = w94 | w115;
assign w514 = w100 | w115;
assign w515 = w98 | w116;
assign w516 = w90 | w116;
assign w517 = w97 | w117;
assign w518 = w100 | w117;
assign w519 = w94 | w118;
assign w520 = w96 | w118;
assign w521 = w98 | w119;
assign w522 = w87 | w119;
assign w523 = w92 | w120;
assign w524 = w99 | w120;
assign w525 = w95 | w121;
assign w526 = w96 | w122;
assign w527 = w100 | w122;
assign w528 = w97 | w123;
assign w529 = w99 | w123;
assign w530 = w94 | w124;
assign w531 = w98 | w124;
assign w532 = w91 | w125;
assign w533 = w95 | w125;
assign w534 = w89 | w126;
assign w535 = ~w127;
assign w536 = ~w128;
assign w537 = w97 | w129;
assign w538 = w93 | w129;
assign w539 = w100 | w129;
assign w540 = w96 | w129;
assign w541 = w94 | w129;
assign w542 = w99 | w129;
assign w543 = w98 | w129;
assign w544 = w127 | w130;
assign w545 = ~w130;
assign w546 = w97 | w131;
assign w547 = w99 | w131;
assign w548 = w96 | w132;
assign w549 = w87 | w132;
assign w550 = w95 | w133;
assign w551 = w93 | w133;
assign w552 = w100 | w134;
assign w553 = w98 | w134;
assign w554 = w75 & w135;
assign w555 = w97 | w136;
assign w556 = w96 | w136;
assign w557 = w99 | w137;
assign w558 = w91 | w137;
assign w559 = w98 | w138;
assign w560 = w94 | w138;
assign w561 = w95 | w139;
assign w562 = w86 | w139;
assign w563 = w179 | w190;
assign w564 = w173 ~| w190;
assign w565 = w175 ~| w190;
assign w566 = w185 | w190;
assign w567 = w184 | w190;
assign w568 = w186 & w192;
assign w569 = w186 ~^ w192;
assign w570 = w171 ~| w193;
assign w571 = w184 | w193;
assign w572 = w183 | w194;
assign w573 = w180 | w194;
assign w574 = w177 ~| w195;
assign w575 = w179 | w196;
assign w576 = w182 | w196;
assign w577 = w191 & w197;
assign w578 = w191 ~^ w197;
assign w579 = w181 | w198;
assign w580 = w180 | w198;
assign w581 = w182 | w199;
assign w582 = w174 | w199;
assign w583 = w179 | w200;
assign w584 = w185 | w200;
assign w585 = w183 | w201;
assign w586 = w175 | w201;
assign w587 = w182 | w202;
assign w588 = w185 | w202;
assign w589 = w179 | w203;
assign w590 = w181 | w203;
assign w591 = w183 | w204;
assign w592 = w172 | w204;
assign w593 = w177 | w205;
assign w594 = w184 | w205;
assign w595 = w180 | w206;
assign w596 = w181 | w207;
assign w597 = w185 | w207;
assign w598 = w182 | w208;
assign w599 = w184 | w208;
assign w600 = w179 | w209;
assign w601 = w183 | w209;
assign w602 = w176 | w210;
assign w603 = w180 | w210;
assign w604 = w174 | w211;
assign w605 = ~w212;
assign w606 = ~w213;
assign w607 = w182 | w214;
assign w608 = w178 | w214;
assign w609 = w185 | w214;
assign w610 = w181 | w214;
assign w611 = w179 | w214;
assign w612 = w184 | w214;
assign w613 = w183 | w214;
assign w614 = w212 | w215;
assign w615 = ~w215;
assign w616 = w182 | w216;
assign w617 = w184 | w216;
assign w618 = w181 | w217;
assign w619 = w172 | w217;
assign w620 = w180 | w218;
assign w621 = w178 | w218;
assign w622 = w185 | w219;
assign w623 = w183 | w219;
assign w624 = w145 & w220;
assign w625 = w182 | w221;
assign w626 = w181 | w221;
assign w627 = w184 | w222;
assign w628 = w176 | w222;
assign w629 = w183 | w223;
assign w630 = w179 | w223;
assign w631 = w180 | w224;
assign w632 = w171 | w224;
assign w633 = w249 | w260;
assign w634 = w243 ~| w260;
assign w635 = w245 ~| w260;
assign w636 = w255 | w260;
assign w637 = w254 | w260;
assign w638 = w256 & w262;
assign w639 = w256 ~^ w262;
assign w640 = w241 ~| w263;
assign w641 = w254 | w263;
assign w642 = w253 | w264;
assign w643 = w250 | w264;
assign w644 = w247 ~| w265;
assign w645 = w249 | w266;
assign w646 = w252 | w266;
assign w647 = w261 & w267;
assign w648 = w261 ~^ w267;
assign w649 = w251 | w268;
assign w650 = w250 | w268;
assign w651 = w252 | w269;
assign w652 = w244 | w269;
assign w653 = w249 | w270;
assign w654 = w255 | w270;
assign w655 = w253 | w271;
assign w656 = w245 | w271;
assign w657 = w252 | w272;
assign w658 = w255 | w272;
assign w659 = w249 | w273;
assign w660 = w251 | w273;
assign w661 = w253 | w274;
assign w662 = w242 | w274;
assign w663 = w247 | w275;
assign w664 = w254 | w275;
assign w665 = w250 | w276;
assign w666 = w251 | w277;
assign w667 = w255 | w277;
assign w668 = w252 | w278;
assign w669 = w254 | w278;
assign w670 = w249 | w279;
assign w671 = w253 | w279;
assign w672 = w246 | w280;
assign w673 = w250 | w280;
assign w674 = w244 | w281;
assign w675 = ~w282;
assign w676 = ~w283;
assign w677 = w252 | w284;
assign w678 = w248 | w284;
assign w679 = w255 | w284;
assign w680 = w251 | w284;
assign w681 = w249 | w284;
assign w682 = w254 | w284;
assign w683 = w253 | w284;
assign w684 = w282 | w285;
assign w685 = ~w285;
assign w686 = w252 | w286;
assign w687 = w254 | w286;
assign w688 = w251 | w287;
assign w689 = w242 | w287;
assign w690 = w250 | w288;
assign w691 = w248 | w288;
assign w692 = w255 | w289;
assign w693 = w253 | w289;
assign w694 = w230 & w290;
assign w695 = w252 | w291;
assign w696 = w251 | w291;
assign w697 = w254 | w292;
assign w698 = w246 | w292;
assign w699 = w253 | w293;
assign w700 = w249 | w293;
assign w701 = w250 | w294;
assign w702 = w241 | w294;
assign w703 = w164 | w299;
assign w704 = w158 ~| w299;
assign w705 = w160 ~| w299;
assign w706 = w170 | w299;
assign w707 = w169 | w299;
assign w708 = w295 & w301;
assign w709 = w295 ~^ w301;
assign w710 = w156 ~| w302;
assign w711 = w169 | w302;
assign w712 = w168 | w303;
assign w713 = w165 | w303;
assign w714 = w162 ~| w304;
assign w715 = w164 | w305;
assign w716 = w167 | w305;
assign w717 = w300 & w306;
assign w718 = w300 ~^ w306;
assign w719 = w166 | w307;
assign w720 = w165 | w307;
assign w721 = w167 | w308;
assign w722 = w159 | w308;
assign w723 = w164 | w309;
assign w724 = w170 | w309;
assign w725 = w168 | w310;
assign w726 = w160 | w310;
assign w727 = w167 | w311;
assign w728 = w170 | w311;
assign w729 = w164 | w312;
assign w730 = w166 | w312;
assign w731 = w168 | w313;
assign w732 = w157 | w313;
assign w733 = w162 | w314;
assign w734 = w169 | w314;
assign w735 = w165 | w315;
assign w736 = w166 | w316;
assign w737 = w170 | w316;
assign w738 = w167 | w317;
assign w739 = w169 | w317;
assign w740 = w164 | w318;
assign w741 = w168 | w318;
assign w742 = w161 | w319;
assign w743 = w165 | w319;
assign w744 = w159 | w320;
assign w745 = ~w321;
assign w746 = ~w322;
assign w747 = w167 | w323;
assign w748 = w163 | w323;
assign w749 = w170 | w323;
assign w750 = w166 | w323;
assign w751 = w164 | w323;
assign w752 = w169 | w323;
assign w753 = w168 | w323;
assign w754 = w321 | w324;
assign w755 = ~w324;
assign w756 = w167 | w325;
assign w757 = w169 | w325;
assign w758 = w166 | w326;
assign w759 = w157 | w326;
assign w760 = w165 | w327;
assign w761 = w163 | w327;
assign w762 = w170 | w328;
assign w763 = w168 | w328;
assign w764 = w167 | w330;
assign w765 = w166 | w330;
assign w766 = w169 | w331;
assign w767 = w161 | w331;
assign w768 = w168 | w332;
assign w769 = w164 | w332;
assign w770 = w165 | w333;
assign w771 = w156 | w333;
assign w772 = w329 & w339;
assign w773 = w377 | w388;
assign w774 = w371 ~| w388;
assign w775 = w373 ~| w388;
assign w776 = w383 | w388;
assign w777 = w382 | w388;
assign w778 = w384 & w390;
assign w779 = w384 ~^ w390;
assign w780 = w369 ~| w391;
assign w781 = w382 | w391;
assign w782 = w381 | w392;
assign w783 = w378 | w392;
assign w784 = w375 ~| w393;
assign w785 = w377 | w394;
assign w786 = w380 | w394;
assign w787 = w389 & w395;
assign w788 = w389 ~^ w395;
assign w789 = w379 | w396;
assign w790 = w378 | w396;
assign w791 = w380 | w397;
assign w792 = w372 | w397;
assign w793 = w377 | w398;
assign w794 = w383 | w398;
assign w795 = w381 | w399;
assign w796 = w373 | w399;
assign w797 = w380 | w400;
assign w798 = w383 | w400;
assign w799 = w377 | w401;
assign w800 = w379 | w401;
assign w801 = w381 | w402;
assign w802 = w370 | w402;
assign w803 = w375 | w403;
assign w804 = w382 | w403;
assign w805 = w378 | w404;
assign w806 = w379 | w405;
assign w807 = w383 | w405;
assign w808 = w380 | w406;
assign w809 = w382 | w406;
assign w810 = w377 | w407;
assign w811 = w381 | w407;
assign w812 = w374 | w408;
assign w813 = w378 | w408;
assign w814 = w372 | w409;
assign w815 = ~w410;
assign w816 = ~w411;
assign w817 = w380 | w412;
assign w818 = w376 | w412;
assign w819 = w383 | w412;
assign w820 = w379 | w412;
assign w821 = w377 | w412;
assign w822 = w382 | w412;
assign w823 = w381 | w412;
assign w824 = w410 | w413;
assign w825 = ~w413;
assign w826 = w380 | w414;
assign w827 = w382 | w414;
assign w828 = w379 | w415;
assign w829 = w370 | w415;
assign w830 = w378 | w416;
assign w831 = w376 | w416;
assign w832 = w383 | w417;
assign w833 = w381 | w417;
assign w834 = w358 & w418;
assign w835 = w380 | w419;
assign w836 = w379 | w419;
assign w837 = w382 | w420;
assign w838 = w374 | w420;
assign w839 = w381 | w421;
assign w840 = w377 | w421;
assign w841 = w378 | w422;
assign w842 = w369 | w422;
assign w843 = w7 & w424;
assign w844 = w0 & w425;
assign w845 = ~w427;
assign w846 = ~w428;
assign w847 = w8 & w430;
assign w848 = w426 ~^ w431;
assign w849 = w427 ~^ w432;
assign w850 = ~w432;
assign w851 = ~w433;
assign w852 = w33 ^ w433;
assign w853 = w7 & w434;
assign w854 = ~w435;
assign w855 = w32 ^ w435;
assign w856 = ~w436;
assign w857 = w34 ^ w436;
assign w858 = ~w437;
assign w859 = w423 ^ w442;
assign w860 = w423 ~| w442;
assign w861 = w431 & w447;
assign w862 = w431 | w447;
assign w863 = w446 ~^ w452;
assign w864 = w446 & w452;
assign w865 = w446 ~| w452;
assign w866 = w444 ~^ w454;
assign w867 = w448 ~^ w459;
assign w868 = w455 ~^ w460;
assign w869 = w455 | w460;
assign w870 = w455 & w460;
assign w871 = w449 ~^ w462;
assign w872 = w449 & w462;
assign w873 = w449 | w462;
assign w874 = w453 ~^ w464;
assign w875 = w453 | w464;
assign w876 = w453 & w464;
assign w877 = w429 ~^ w466;
assign w878 = w454 | w467;
assign w879 = w454 & w467;
assign w880 = w458 ~^ w470;
assign w881 = w458 & w470;
assign w882 = w458 | w470;
assign w883 = w441 ~^ w471;
assign w884 = w457 ~^ w472;
assign w885 = w465 ~^ w475;
assign w886 = w465 ~| w475;
assign w887 = w459 & w476;
assign w888 = w459 | w476;
assign w889 = w469 ~^ w477;
assign w890 = w461 ~^ w478;
assign w891 = w468 ~^ w479;
assign w892 = w468 & w479;
assign w893 = w468 | w479;
assign w894 = w471 | w481;
assign w895 = w471 & w481;
assign w896 = w472 | w485;
assign w897 = w472 & w485;
assign w898 = w473 ~^ w486;
assign w899 = w473 | w486;
assign w900 = w473 & w486;
assign w901 = w482 ~^ w487;
assign w902 = w482 & w487;
assign w903 = w482 ~| w487;
assign w904 = w456 ~^ w488;
assign w905 = w456 | w488;
assign w906 = w456 & w488;
assign w907 = w477 & w489;
assign w908 = w477 | w489;
assign w909 = w480 ~^ w490;
assign w910 = w480 & w490;
assign w911 = w480 | w490;
assign w912 = w478 | w491;
assign w913 = w478 & w491;
assign w914 = w450 ~^ w492;
assign w915 = w463 & w492;
assign w916 = w463 | w492;
assign w917 = w77 & w494;
assign w918 = w70 & w495;
assign w919 = ~w497;
assign w920 = ~w498;
assign w921 = w78 & w500;
assign w922 = w496 ~^ w501;
assign w923 = w497 ~^ w502;
assign w924 = ~w502;
assign w925 = ~w503;
assign w926 = w103 ^ w503;
assign w927 = w77 & w504;
assign w928 = ~w505;
assign w929 = w102 ^ w505;
assign w930 = ~w506;
assign w931 = w104 ^ w506;
assign w932 = ~w507;
assign w933 = w493 ^ w512;
assign w934 = w493 ~| w512;
assign w935 = w501 & w517;
assign w936 = w501 | w517;
assign w937 = w516 ~^ w522;
assign w938 = w516 & w522;
assign w939 = w516 ~| w522;
assign w940 = w514 ~^ w524;
assign w941 = w518 ~^ w529;
assign w942 = w525 ~^ w530;
assign w943 = w525 | w530;
assign w944 = w525 & w530;
assign w945 = w519 ~^ w532;
assign w946 = w519 & w532;
assign w947 = w519 | w532;
assign w948 = w523 ~^ w534;
assign w949 = w523 | w534;
assign w950 = w523 & w534;
assign w951 = w499 ~^ w536;
assign w952 = w524 | w537;
assign w953 = w524 & w537;
assign w954 = w528 ~^ w540;
assign w955 = w528 & w540;
assign w956 = w528 | w540;
assign w957 = w511 ~^ w541;
assign w958 = w527 ~^ w542;
assign w959 = w535 ~^ w545;
assign w960 = w535 ~| w545;
assign w961 = w529 & w546;
assign w962 = w529 | w546;
assign w963 = w539 ~^ w547;
assign w964 = w531 ~^ w548;
assign w965 = w538 ~^ w549;
assign w966 = w538 & w549;
assign w967 = w538 | w549;
assign w968 = w541 | w551;
assign w969 = w541 & w551;
assign w970 = w542 | w555;
assign w971 = w542 & w555;
assign w972 = w543 ~^ w556;
assign w973 = w543 | w556;
assign w974 = w543 & w556;
assign w975 = w552 ~^ w557;
assign w976 = w552 & w557;
assign w977 = w552 ~| w557;
assign w978 = w526 ~^ w558;
assign w979 = w526 | w558;
assign w980 = w526 & w558;
assign w981 = w547 & w559;
assign w982 = w547 | w559;
assign w983 = w550 ~^ w560;
assign w984 = w550 & w560;
assign w985 = w550 | w560;
assign w986 = w548 | w561;
assign w987 = w548 & w561;
assign w988 = w520 ~^ w562;
assign w989 = w533 & w562;
assign w990 = w533 | w562;
assign w991 = w147 & w564;
assign w992 = w140 & w565;
assign w993 = ~w567;
assign w994 = ~w568;
assign w995 = w148 & w570;
assign w996 = w566 ~^ w571;
assign w997 = w567 ~^ w572;
assign w998 = ~w572;
assign w999 = ~w573;
assign w1000 = w188 ^ w573;
assign w1001 = w147 & w574;
assign w1002 = ~w575;
assign w1003 = w187 ^ w575;
assign w1004 = ~w576;
assign w1005 = w189 ^ w576;
assign w1006 = ~w577;
assign w1007 = w563 ^ w582;
assign w1008 = w563 ~| w582;
assign w1009 = w571 & w587;
assign w1010 = w571 | w587;
assign w1011 = w586 ~^ w592;
assign w1012 = w586 & w592;
assign w1013 = w586 ~| w592;
assign w1014 = w584 ~^ w594;
assign w1015 = w588 ~^ w599;
assign w1016 = w595 ~^ w600;
assign w1017 = w595 | w600;
assign w1018 = w595 & w600;
assign w1019 = w589 ~^ w602;
assign w1020 = w589 & w602;
assign w1021 = w589 | w602;
assign w1022 = w593 ~^ w604;
assign w1023 = w593 | w604;
assign w1024 = w593 & w604;
assign w1025 = w569 ~^ w606;
assign w1026 = w594 | w607;
assign w1027 = w594 & w607;
assign w1028 = w598 ~^ w610;
assign w1029 = w598 & w610;
assign w1030 = w598 | w610;
assign w1031 = w581 ~^ w611;
assign w1032 = w597 ~^ w612;
assign w1033 = w605 ~^ w615;
assign w1034 = w605 ~| w615;
assign w1035 = w599 & w616;
assign w1036 = w599 | w616;
assign w1037 = w609 ~^ w617;
assign w1038 = w601 ~^ w618;
assign w1039 = w608 ~^ w619;
assign w1040 = w608 & w619;
assign w1041 = w608 | w619;
assign w1042 = w611 | w621;
assign w1043 = w611 & w621;
assign w1044 = w554 ~^ w624;
assign w1045 = w612 | w625;
assign w1046 = w612 & w625;
assign w1047 = w613 ~^ w626;
assign w1048 = w613 | w626;
assign w1049 = w613 & w626;
assign w1050 = w622 ~^ w627;
assign w1051 = w622 & w627;
assign w1052 = w622 ~| w627;
assign w1053 = w596 ~^ w628;
assign w1054 = w596 | w628;
assign w1055 = w596 & w628;
assign w1056 = w617 & w629;
assign w1057 = w617 | w629;
assign w1058 = w620 ~^ w630;
assign w1059 = w620 & w630;
assign w1060 = w620 | w630;
assign w1061 = w618 | w631;
assign w1062 = w618 & w631;
assign w1063 = w590 ~^ w632;
assign w1064 = w603 & w632;
assign w1065 = w603 | w632;
assign w1066 = w232 & w634;
assign w1067 = w225 & w635;
assign w1068 = ~w637;
assign w1069 = ~w638;
assign w1070 = w233 & w640;
assign w1071 = w636 ~^ w641;
assign w1072 = w637 ~^ w642;
assign w1073 = ~w642;
assign w1074 = ~w643;
assign w1075 = w258 ^ w643;
assign w1076 = w232 & w644;
assign w1077 = ~w645;
assign w1078 = w257 ^ w645;
assign w1079 = ~w646;
assign w1080 = w259 ^ w646;
assign w1081 = ~w647;
assign w1082 = w633 ^ w652;
assign w1083 = w633 ~| w652;
assign w1084 = w641 & w657;
assign w1085 = w641 | w657;
assign w1086 = w656 ~^ w662;
assign w1087 = w656 & w662;
assign w1088 = w656 ~| w662;
assign w1089 = w654 ~^ w664;
assign w1090 = w658 ~^ w669;
assign w1091 = w665 ~^ w670;
assign w1092 = w665 | w670;
assign w1093 = w665 & w670;
assign w1094 = w659 ~^ w672;
assign w1095 = w659 & w672;
assign w1096 = w659 | w672;
assign w1097 = w663 ~^ w674;
assign w1098 = w663 | w674;
assign w1099 = w663 & w674;
assign w1100 = w639 ~^ w676;
assign w1101 = w664 | w677;
assign w1102 = w664 & w677;
assign w1103 = w668 ~^ w680;
assign w1104 = w668 & w680;
assign w1105 = w668 | w680;
assign w1106 = w651 ~^ w681;
assign w1107 = w667 ~^ w682;
assign w1108 = w675 ~^ w685;
assign w1109 = w675 ~| w685;
assign w1110 = w669 & w686;
assign w1111 = w669 | w686;
assign w1112 = w679 ~^ w687;
assign w1113 = w671 ~^ w688;
assign w1114 = w678 ~^ w689;
assign w1115 = w678 & w689;
assign w1116 = w678 | w689;
assign w1117 = w681 | w691;
assign w1118 = w681 & w691;
assign w1119 = ~w694;
assign w1120 = w682 | w695;
assign w1121 = w682 & w695;
assign w1122 = w683 ~^ w696;
assign w1123 = w683 | w696;
assign w1124 = w683 & w696;
assign w1125 = w692 ~^ w697;
assign w1126 = w692 & w697;
assign w1127 = w692 ~| w697;
assign w1128 = w666 ~^ w698;
assign w1129 = w666 | w698;
assign w1130 = w666 & w698;
assign w1131 = w687 & w699;
assign w1132 = w687 | w699;
assign w1133 = w690 ~^ w700;
assign w1134 = w690 & w700;
assign w1135 = w690 | w700;
assign w1136 = w688 | w701;
assign w1137 = w688 & w701;
assign w1138 = w660 ~^ w702;
assign w1139 = w673 & w702;
assign w1140 = w673 | w702;
assign w1141 = w341 & w704;
assign w1142 = w334 & w705;
assign w1143 = ~w707;
assign w1144 = ~w708;
assign w1145 = w342 & w710;
assign w1146 = w706 ~^ w711;
assign w1147 = w707 ~^ w712;
assign w1148 = ~w712;
assign w1149 = ~w713;
assign w1150 = w297 ^ w713;
assign w1151 = w341 & w714;
assign w1152 = ~w715;
assign w1153 = w296 ^ w715;
assign w1154 = ~w716;
assign w1155 = w298 ^ w716;
assign w1156 = ~w717;
assign w1157 = w703 ^ w722;
assign w1158 = w703 ~| w722;
assign w1159 = w711 & w727;
assign w1160 = w711 | w727;
assign w1161 = w726 ~^ w732;
assign w1162 = w726 & w732;
assign w1163 = w726 ~| w732;
assign w1164 = w724 ~^ w734;
assign w1165 = w728 ~^ w739;
assign w1166 = w735 ~^ w740;
assign w1167 = w735 | w740;
assign w1168 = w735 & w740;
assign w1169 = w729 ~^ w742;
assign w1170 = w729 & w742;
assign w1171 = w729 | w742;
assign w1172 = w733 ~^ w744;
assign w1173 = w733 | w744;
assign w1174 = w733 & w744;
assign w1175 = w709 ~^ w746;
assign w1176 = w734 | w747;
assign w1177 = w734 & w747;
assign w1178 = w738 ~^ w750;
assign w1179 = w738 & w750;
assign w1180 = w738 | w750;
assign w1181 = w721 ~^ w751;
assign w1182 = w737 ~^ w752;
assign w1183 = w745 ~^ w755;
assign w1184 = w745 ~| w755;
assign w1185 = w739 & w756;
assign w1186 = w739 | w756;
assign w1187 = w749 ~^ w757;
assign w1188 = w741 ~^ w758;
assign w1189 = w748 ~^ w759;
assign w1190 = w748 & w759;
assign w1191 = w748 | w759;
assign w1192 = w751 | w761;
assign w1193 = w751 & w761;
assign w1194 = w752 | w764;
assign w1195 = w752 & w764;
assign w1196 = w753 ~^ w765;
assign w1197 = w753 | w765;
assign w1198 = w753 & w765;
assign w1199 = w762 ~^ w766;
assign w1200 = w762 & w766;
assign w1201 = w762 ~| w766;
assign w1202 = w736 ~^ w767;
assign w1203 = w736 | w767;
assign w1204 = w736 & w767;
assign w1205 = w757 & w768;
assign w1206 = w757 | w768;
assign w1207 = w760 ~^ w769;
assign w1208 = w760 & w769;
assign w1209 = w760 | w769;
assign w1210 = w758 | w770;
assign w1211 = w758 & w770;
assign w1212 = w730 ~^ w771;
assign w1213 = w743 & w771;
assign w1214 = w743 | w771;
assign w1215 = w694 ~^ w772;
assign w1216 = ~w772;
assign w1217 = w360 & w774;
assign w1218 = w353 & w775;
assign w1219 = ~w777;
assign w1220 = ~w778;
assign w1221 = w361 & w780;
assign w1222 = w776 ~^ w781;
assign w1223 = w777 ~^ w782;
assign w1224 = ~w782;
assign w1225 = ~w783;
assign w1226 = w386 ^ w783;
assign w1227 = w360 & w784;
assign w1228 = ~w785;
assign w1229 = w385 ^ w785;
assign w1230 = ~w786;
assign w1231 = w387 ^ w786;
assign w1232 = ~w787;
assign w1233 = w773 ^ w792;
assign w1234 = w773 ~| w792;
assign w1235 = w781 & w797;
assign w1236 = w781 | w797;
assign w1237 = w796 ~^ w802;
assign w1238 = w796 & w802;
assign w1239 = w796 ~| w802;
assign w1240 = w794 ~^ w804;
assign w1241 = w798 ~^ w809;
assign w1242 = w805 ~^ w810;
assign w1243 = w805 | w810;
assign w1244 = w805 & w810;
assign w1245 = w799 ~^ w812;
assign w1246 = w799 & w812;
assign w1247 = w799 | w812;
assign w1248 = w803 ~^ w814;
assign w1249 = w803 | w814;
assign w1250 = w803 & w814;
assign w1251 = w779 ~^ w816;
assign w1252 = w804 | w817;
assign w1253 = w804 & w817;
assign w1254 = w808 ~^ w820;
assign w1255 = w808 & w820;
assign w1256 = w808 | w820;
assign w1257 = w791 ~^ w821;
assign w1258 = w807 ~^ w822;
assign w1259 = w815 ~^ w825;
assign w1260 = w815 ~| w825;
assign w1261 = w809 & w826;
assign w1262 = w809 | w826;
assign w1263 = w819 ~^ w827;
assign w1264 = w811 ~^ w828;
assign w1265 = w818 ~^ w829;
assign w1266 = w818 & w829;
assign w1267 = w818 | w829;
assign w1268 = w821 | w831;
assign w1269 = w821 & w831;
assign w1270 = w554 & w834;
assign w1271 = w554 | w834;
assign w1272 = w822 | w835;
assign w1273 = w822 & w835;
assign w1274 = w823 ~^ w836;
assign w1275 = w823 | w836;
assign w1276 = w823 & w836;
assign w1277 = w832 ~^ w837;
assign w1278 = w832 & w837;
assign w1279 = w832 ~| w837;
assign w1280 = w806 ~^ w838;
assign w1281 = w806 | w838;
assign w1282 = w806 & w838;
assign w1283 = w827 & w839;
assign w1284 = w827 | w839;
assign w1285 = w830 ~^ w840;
assign w1286 = w830 & w840;
assign w1287 = w830 | w840;
assign w1288 = w828 | w841;
assign w1289 = w828 & w841;
assign w1290 = w800 ~^ w842;
assign w1291 = w813 & w842;
assign w1292 = w813 | w842;
assign w1293 = in5[0] ~^ w843;
assign w1294 = w843 & in5[0];
assign w1295 = in5[1] ~| w844;
assign w1296 = ~w844;
assign w1297 = w447 ~^ w848;
assign w1298 = ~w849;
assign w1299 = w845 & w850;
assign w1300 = w33 & w851;
assign w1301 = w32 & w854;
assign w1302 = w34 & w856;
assign w1303 = w15 & w859;
assign w1304 = w6 & w860;
assign w1305 = w426 | w861;
assign w1306 = w855 ^ w863;
assign w1307 = w855 ~| w864;
assign w1308 = w467 ~^ w866;
assign w1309 = w476 ~^ w867;
assign w1310 = w439 ~^ w868;
assign w1311 = w439 | w870;
assign w1312 = w440 ~^ w871;
assign w1313 = w440 | w872;
assign w1314 = w443 ~^ w874;
assign w1315 = w443 | w876;
assign w1316 = w444 | w879;
assign w1317 = w451 ~^ w880;
assign w1318 = w451 | w881;
assign w1319 = w481 ~^ w883;
assign w1320 = w485 ~^ w884;
assign w1321 = w448 | w887;
assign w1322 = w489 ~^ w889;
assign w1323 = w491 ~^ w890;
assign w1324 = w428 ~^ w891;
assign w1325 = w846 | w892;
assign w1326 = w441 | w895;
assign w1327 = w457 | w897;
assign w1328 = w445 ~^ w904;
assign w1329 = w445 | w906;
assign w1330 = w469 | w907;
assign w1331 = w438 ~^ w909;
assign w1332 = w438 | w910;
assign w1333 = w461 | w913;
assign w1334 = w463 ~^ w914;
assign w1335 = w450 | w915;
assign w1336 = ~w917;
assign w1337 = w517 ~^ w922;
assign w1338 = ~w923;
assign w1339 = w919 & w924;
assign w1340 = w103 & w925;
assign w1341 = w102 & w928;
assign w1342 = w104 & w930;
assign w1343 = w85 & w933;
assign w1344 = w76 & w934;
assign w1345 = w496 | w935;
assign w1346 = w929 ^ w937;
assign w1347 = w929 ~| w938;
assign w1348 = w537 ~^ w940;
assign w1349 = w546 ~^ w941;
assign w1350 = w509 ~^ w942;
assign w1351 = w509 | w944;
assign w1352 = w510 ~^ w945;
assign w1353 = w510 | w946;
assign w1354 = w513 ~^ w948;
assign w1355 = w513 | w950;
assign w1356 = w514 | w953;
assign w1357 = w521 ~^ w954;
assign w1358 = w521 | w955;
assign w1359 = w551 ~^ w957;
assign w1360 = w555 ~^ w958;
assign w1361 = w518 | w961;
assign w1362 = w559 ~^ w963;
assign w1363 = w561 ~^ w964;
assign w1364 = w498 ~^ w965;
assign w1365 = w920 | w966;
assign w1366 = w511 | w969;
assign w1367 = w527 | w971;
assign w1368 = w515 ~^ w978;
assign w1369 = w515 | w980;
assign w1370 = w539 | w981;
assign w1371 = w508 ~^ w983;
assign w1372 = w508 | w984;
assign w1373 = w531 | w987;
assign w1374 = w533 ~^ w988;
assign w1375 = w520 | w989;
assign w1376 = w917 ~| w991;
assign w1377 = ~w991;
assign w1378 = w918 ~^ w992;
assign w1379 = w918 & w992;
assign w1380 = w918 | w992;
assign w1381 = w587 ~^ w996;
assign w1382 = ~w997;
assign w1383 = w993 & w998;
assign w1384 = w188 & w999;
assign w1385 = w187 & w1002;
assign w1386 = w189 & w1004;
assign w1387 = w155 & w1007;
assign w1388 = w146 & w1008;
assign w1389 = w566 | w1009;
assign w1390 = w1003 ^ w1011;
assign w1391 = w1003 ~| w1012;
assign w1392 = w607 ~^ w1014;
assign w1393 = w616 ~^ w1015;
assign w1394 = w579 ~^ w1016;
assign w1395 = w579 | w1018;
assign w1396 = w580 ~^ w1019;
assign w1397 = w580 | w1020;
assign w1398 = w583 ~^ w1022;
assign w1399 = w583 | w1024;
assign w1400 = w584 | w1027;
assign w1401 = w591 ~^ w1028;
assign w1402 = w591 | w1029;
assign w1403 = w621 ~^ w1031;
assign w1404 = w625 ~^ w1032;
assign w1405 = w588 | w1035;
assign w1406 = w629 ~^ w1037;
assign w1407 = w631 ~^ w1038;
assign w1408 = w568 ~^ w1039;
assign w1409 = w994 | w1040;
assign w1410 = w581 | w1043;
assign w1411 = w834 ~^ w1044;
assign w1412 = w597 | w1046;
assign w1413 = w585 ~^ w1053;
assign w1414 = w585 | w1055;
assign w1415 = w609 | w1056;
assign w1416 = w578 ~^ w1058;
assign w1417 = w578 | w1059;
assign w1418 = w601 | w1062;
assign w1419 = w603 ~^ w1063;
assign w1420 = w590 | w1064;
assign w1421 = w1067 ~^ in5[1];
assign w1422 = ~w1067;
assign w1423 = w657 ~^ w1071;
assign w1424 = ~w1072;
assign w1425 = w1068 & w1073;
assign w1426 = w258 & w1074;
assign w1427 = w1076 ~^ in5[2];
assign w1428 = ~w1076;
assign w1429 = w257 & w1077;
assign w1430 = w259 & w1079;
assign w1431 = w240 & w1082;
assign w1432 = w231 & w1083;
assign w1433 = w636 | w1084;
assign w1434 = w1078 ^ w1086;
assign w1435 = w1078 ~| w1087;
assign w1436 = w677 ~^ w1089;
assign w1437 = w686 ~^ w1090;
assign w1438 = w649 ~^ w1091;
assign w1439 = w649 | w1093;
assign w1440 = w650 ~^ w1094;
assign w1441 = w650 | w1095;
assign w1442 = w653 ~^ w1097;
assign w1443 = w653 | w1099;
assign w1444 = w654 | w1102;
assign w1445 = w661 ~^ w1103;
assign w1446 = w661 | w1104;
assign w1447 = w691 ~^ w1106;
assign w1448 = w695 ~^ w1107;
assign w1449 = w658 | w1110;
assign w1450 = w699 ~^ w1112;
assign w1451 = w701 ~^ w1113;
assign w1452 = w638 ~^ w1114;
assign w1453 = w1069 | w1115;
assign w1454 = w651 | w1118;
assign w1455 = w667 | w1121;
assign w1456 = w655 ~^ w1128;
assign w1457 = w655 | w1130;
assign w1458 = w679 | w1131;
assign w1459 = w648 ~^ w1133;
assign w1460 = w648 | w1134;
assign w1461 = w671 | w1137;
assign w1462 = w673 ~^ w1138;
assign w1463 = w660 | w1139;
assign w1464 = w1066 & w1141;
assign w1465 = ~w1141;
assign w1466 = w727 ~^ w1146;
assign w1467 = ~w1147;
assign w1468 = w1143 & w1148;
assign w1469 = w297 & w1149;
assign w1470 = w296 & w1152;
assign w1471 = w298 & w1154;
assign w1472 = w349 & w1157;
assign w1473 = w340 & w1158;
assign w1474 = w706 | w1159;
assign w1475 = w1153 ^ w1161;
assign w1476 = w1153 ~| w1162;
assign w1477 = w747 ~^ w1164;
assign w1478 = w756 ~^ w1165;
assign w1479 = w719 ~^ w1166;
assign w1480 = w719 | w1168;
assign w1481 = w720 ~^ w1169;
assign w1482 = w720 | w1170;
assign w1483 = w723 ~^ w1172;
assign w1484 = w723 | w1174;
assign w1485 = w724 | w1177;
assign w1486 = w731 ~^ w1178;
assign w1487 = w731 | w1179;
assign w1488 = w761 ~^ w1181;
assign w1489 = w764 ~^ w1182;
assign w1490 = w728 | w1185;
assign w1491 = w768 ~^ w1187;
assign w1492 = w770 ~^ w1188;
assign w1493 = w708 ~^ w1189;
assign w1494 = w1144 | w1190;
assign w1495 = w721 | w1193;
assign w1496 = w737 | w1195;
assign w1497 = w725 ~^ w1202;
assign w1498 = w725 | w1204;
assign w1499 = w749 | w1205;
assign w1500 = w718 ~^ w1207;
assign w1501 = w718 | w1208;
assign w1502 = w741 | w1211;
assign w1503 = w743 ~^ w1212;
assign w1504 = w730 | w1213;
assign w1505 = w484 ~^ w1215;
assign w1506 = w1119 | w1216;
assign w1507 = w991 ~^ w1217;
assign w1508 = ~w1217;
assign w1509 = w1142 ~^ w1218;
assign w1510 = w1142 | w1218;
assign w1511 = w1142 & w1218;
assign w1512 = w995 ~^ w1221;
assign w1513 = w847 & w1221;
assign w1514 = w847 | w1221;
assign w1515 = w797 ~^ w1222;
assign w1516 = ~w1223;
assign w1517 = w1219 & w1224;
assign w1518 = w386 & w1225;
assign w1519 = w385 & w1228;
assign w1520 = w387 & w1230;
assign w1521 = w368 & w1233;
assign w1522 = w359 & w1234;
assign w1523 = w776 | w1235;
assign w1524 = w1229 ^ w1237;
assign w1525 = w1229 ~| w1238;
assign w1526 = w817 ~^ w1240;
assign w1527 = w826 ~^ w1241;
assign w1528 = w789 ~^ w1242;
assign w1529 = w789 | w1244;
assign w1530 = w790 ~^ w1245;
assign w1531 = w790 | w1246;
assign w1532 = w793 ~^ w1248;
assign w1533 = w793 | w1250;
assign w1534 = w794 | w1253;
assign w1535 = w801 ~^ w1254;
assign w1536 = w801 | w1255;
assign w1537 = w831 ~^ w1257;
assign w1538 = w835 ~^ w1258;
assign w1539 = w798 | w1261;
assign w1540 = w839 ~^ w1263;
assign w1541 = w841 ~^ w1264;
assign w1542 = w778 ~^ w1265;
assign w1543 = w1220 | w1266;
assign w1544 = w791 | w1269;
assign w1545 = w624 & w1271;
assign w1546 = w807 | w1273;
assign w1547 = w795 ~^ w1280;
assign w1548 = w795 | w1282;
assign w1549 = w819 | w1283;
assign w1550 = w788 ~^ w1285;
assign w1551 = w788 | w1286;
assign w1552 = w811 | w1289;
assign w1553 = w813 ~^ w1290;
assign w1554 = w800 | w1291;
assign w1555 = ~w1293;
assign w1556 = w1070 ~^ w1294;
assign w1557 = ~w1294;
assign w1558 = w350 | w1296;
assign w1559 = w885 ~^ w1299;
assign w1560 = w474 & w1299;
assign w1561 = w877 ~^ w1300;
assign w1562 = w58 ~| w1300;
assign w1563 = ~w1300;
assign w1564 = w852 ~^ w1301;
assign w1565 = ~w1301;
assign w1566 = w849 ~^ w1302;
assign w1567 = w1298 ~| w1302;
assign w1568 = ~w1302;
assign w1569 = w927 ~^ w1303;
assign w1570 = w927 & w1303;
assign w1571 = w927 ~| w1303;
assign w1572 = w862 & w1305;
assign w1573 = w14 & w1306;
assign w1574 = w865 | w1307;
assign w1575 = ~w1308;
assign w1576 = w869 & w1311;
assign w1577 = ~w1312;
assign w1578 = w873 & w1313;
assign w1579 = w875 & w1315;
assign w1580 = w878 & w1316;
assign w1581 = w882 & w1318;
assign w1582 = w888 & w1321;
assign w1583 = ~w1324;
assign w1584 = w893 & w1325;
assign w1585 = w894 & w1326;
assign w1586 = w896 & w1327;
assign w1587 = ~w1328;
assign w1588 = w905 & w1329;
assign w1589 = w908 & w1330;
assign w1590 = ~w1331;
assign w1591 = w911 & w1332;
assign w1592 = w912 & w1333;
assign w1593 = w1319 ~^ w1334;
assign w1594 = w1319 ~| w1334;
assign w1595 = w1319 & w1334;
assign w1596 = w916 & w1335;
assign w1597 = w959 ~^ w1339;
assign w1598 = w544 & w1339;
assign w1599 = w951 ~^ w1340;
assign w1600 = w128 ~| w1340;
assign w1601 = ~w1340;
assign w1602 = w926 ~^ w1341;
assign w1603 = ~w1341;
assign w1604 = w923 ~^ w1342;
assign w1605 = w1338 ~| w1342;
assign w1606 = ~w1342;
assign w1607 = w936 & w1345;
assign w1608 = w84 & w1346;
assign w1609 = w939 | w1347;
assign w1610 = ~w1348;
assign w1611 = w943 & w1351;
assign w1612 = ~w1352;
assign w1613 = w947 & w1353;
assign w1614 = w949 & w1355;
assign w1615 = w952 & w1356;
assign w1616 = w956 & w1358;
assign w1617 = w962 & w1361;
assign w1618 = ~w1364;
assign w1619 = w967 & w1365;
assign w1620 = w968 & w1366;
assign w1621 = w970 & w1367;
assign w1622 = ~w1368;
assign w1623 = w979 & w1369;
assign w1624 = w982 & w1370;
assign w1625 = ~w1371;
assign w1626 = w985 & w1372;
assign w1627 = w986 & w1373;
assign w1628 = w1359 ~^ w1374;
assign w1629 = w1359 ~| w1374;
assign w1630 = w1359 & w1374;
assign w1631 = w990 & w1375;
assign w1632 = w1336 | w1377;
assign w1633 = w921 ~^ w1378;
assign w1634 = w921 & w1380;
assign w1635 = w1033 ~^ w1383;
assign w1636 = w614 & w1383;
assign w1637 = w1025 ~^ w1384;
assign w1638 = w213 ~| w1384;
assign w1639 = ~w1384;
assign w1640 = w1000 ~^ w1385;
assign w1641 = ~w1385;
assign w1642 = w997 ~^ w1386;
assign w1643 = w1382 ~| w1386;
assign w1644 = ~w1386;
assign w1645 = w853 ~^ w1387;
assign w1646 = w853 | w1387;
assign w1647 = w853 & w1387;
assign w1648 = w1010 & w1389;
assign w1649 = w154 & w1390;
assign w1650 = w1013 | w1391;
assign w1651 = ~w1392;
assign w1652 = w1017 & w1395;
assign w1653 = ~w1396;
assign w1654 = w1021 & w1397;
assign w1655 = w1023 & w1399;
assign w1656 = w1026 & w1400;
assign w1657 = w1030 & w1402;
assign w1658 = w1036 & w1405;
assign w1659 = ~w1408;
assign w1660 = w1041 & w1409;
assign w1661 = w1042 & w1410;
assign w1662 = w1045 & w1412;
assign w1663 = ~w1413;
assign w1664 = w1054 & w1414;
assign w1665 = w1057 & w1415;
assign w1666 = ~w1416;
assign w1667 = w1060 & w1417;
assign w1668 = w1061 & w1418;
assign w1669 = w1403 ~^ w1419;
assign w1670 = w1403 ~| w1419;
assign w1671 = w1403 & w1419;
assign w1672 = w1065 & w1420;
assign w1673 = w844 ^ w1421;
assign w1674 = w1295 | w1422;
assign w1675 = w1108 ~^ w1425;
assign w1676 = w684 & w1425;
assign w1677 = w1100 ~^ w1426;
assign w1678 = w283 ~| w1426;
assign w1679 = ~w1426;
assign w1680 = w351 | w1428;
assign w1681 = w1075 ~^ w1429;
assign w1682 = ~w1429;
assign w1683 = w1072 ~^ w1430;
assign w1684 = w1424 ~| w1430;
assign w1685 = ~w1430;
assign w1686 = w1343 ~^ w1431;
assign w1687 = w1343 & w1431;
assign w1688 = w1343 | w1431;
assign w1689 = w1432 ~^ in5[3];
assign w1690 = ~w1432;
assign w1691 = w1085 & w1433;
assign w1692 = w239 & w1434;
assign w1693 = w1088 | w1435;
assign w1694 = ~w1436;
assign w1695 = w1092 & w1439;
assign w1696 = ~w1440;
assign w1697 = w1096 & w1441;
assign w1698 = w1098 & w1443;
assign w1699 = w1101 & w1444;
assign w1700 = w1105 & w1446;
assign w1701 = w1111 & w1449;
assign w1702 = ~w1452;
assign w1703 = w1116 & w1453;
assign w1704 = w1117 & w1454;
assign w1705 = w1120 & w1455;
assign w1706 = ~w1456;
assign w1707 = w1129 & w1457;
assign w1708 = w1132 & w1458;
assign w1709 = ~w1459;
assign w1710 = w1135 & w1460;
assign w1711 = w1136 & w1461;
assign w1712 = w1447 ~^ w1462;
assign w1713 = w1447 ~| w1462;
assign w1714 = w1447 & w1462;
assign w1715 = w1140 & w1463;
assign w1716 = w1066 ~^ w1465;
assign w1717 = w1183 ~^ w1468;
assign w1718 = w754 & w1468;
assign w1719 = w1175 ~^ w1469;
assign w1720 = w322 ~| w1469;
assign w1721 = ~w1469;
assign w1722 = w1150 ~^ w1470;
assign w1723 = ~w1470;
assign w1724 = w1147 ~^ w1471;
assign w1725 = w1467 ~| w1471;
assign w1726 = ~w1471;
assign w1727 = w1227 ~^ w1472;
assign w1728 = w1227 | w1472;
assign w1729 = w1227 & w1472;
assign w1730 = w1388 ~^ w1473;
assign w1731 = w1388 | w1473;
assign w1732 = w1388 & w1473;
assign w1733 = w1160 & w1474;
assign w1734 = w348 & w1475;
assign w1735 = w1163 | w1476;
assign w1736 = ~w1477;
assign w1737 = w1167 & w1480;
assign w1738 = ~w1481;
assign w1739 = w1171 & w1482;
assign w1740 = w1173 & w1484;
assign w1741 = w1176 & w1485;
assign w1742 = w1180 & w1487;
assign w1743 = w1186 & w1490;
assign w1744 = ~w1493;
assign w1745 = w1191 & w1494;
assign w1746 = w1192 & w1495;
assign w1747 = w1194 & w1496;
assign w1748 = ~w1497;
assign w1749 = w1203 & w1498;
assign w1750 = w1206 & w1499;
assign w1751 = ~w1500;
assign w1752 = w1209 & w1501;
assign w1753 = w1210 & w1502;
assign w1754 = w1488 ~^ w1503;
assign w1755 = w1488 ~| w1503;
assign w1756 = w1488 & w1503;
assign w1757 = w1214 & w1504;
assign w1758 = ~w1506;
assign w1759 = w917 ~^ w1507;
assign w1760 = w1376 | w1508;
assign w1761 = w1145 ~^ w1509;
assign w1762 = w1145 & w1510;
assign w1763 = w847 ~^ w1512;
assign w1764 = w995 & w1514;
assign w1765 = w1259 ~^ w1517;
assign w1766 = w824 & w1517;
assign w1767 = w1251 ~^ w1518;
assign w1768 = w411 ~| w1518;
assign w1769 = ~w1518;
assign w1770 = w1226 ~^ w1519;
assign w1771 = ~w1519;
assign w1772 = w1223 ~^ w1520;
assign w1773 = w1516 ~| w1520;
assign w1774 = ~w1520;
assign w1775 = w1304 ~^ w1522;
assign w1776 = w1304 & w1522;
assign w1777 = w1304 | w1522;
assign w1778 = w1236 & w1523;
assign w1779 = w367 & w1524;
assign w1780 = w1239 | w1525;
assign w1781 = ~w1526;
assign w1782 = w1243 & w1529;
assign w1783 = ~w1530;
assign w1784 = w1247 & w1531;
assign w1785 = w1249 & w1533;
assign w1786 = w1252 & w1534;
assign w1787 = w1256 & w1536;
assign w1788 = w1262 & w1539;
assign w1789 = ~w1542;
assign w1790 = w1267 & w1543;
assign w1791 = w1268 & w1544;
assign w1792 = w1270 | w1545;
assign w1793 = w1272 & w1546;
assign w1794 = ~w1547;
assign w1795 = w1281 & w1548;
assign w1796 = w1284 & w1549;
assign w1797 = ~w1550;
assign w1798 = w1287 & w1551;
assign w1799 = w1288 & w1552;
assign w1800 = w1537 ~^ w1553;
assign w1801 = w1537 ~| w1553;
assign w1802 = w1537 & w1553;
assign w1803 = w1292 & w1554;
assign w1804 = w1328 ~^ w1559;
assign w1805 = ~w1559;
assign w1806 = w886 | w1560;
assign w1807 = w429 | w1562;
assign w1808 = w466 | w1563;
assign w1809 = w1314 ~^ w1564;
assign w1810 = w852 & w1565;
assign w1811 = w852 ~| w1565;
assign w1812 = w849 | w1568;
assign w1813 = w1427 ~^ w1569;
assign w1814 = w1427 ~| w1571;
assign w1815 = ~w1573;
assign w1816 = w2 & w1574;
assign w1817 = w1566 ~^ w1576;
assign w1818 = w1567 | w1576;
assign w1819 = w857 ~^ w1578;
assign w1820 = w857 | w1578;
assign w1821 = w857 & w1578;
assign w1822 = w1312 ~^ w1579;
assign w1823 = w1312 ~| w1579;
assign w1824 = ~w1579;
assign w1825 = w1309 ~^ w1580;
assign w1826 = w437 ~^ w1581;
assign w1827 = w858 | w1581;
assign w1828 = ~w1581;
assign w1829 = w483 ~^ w1582;
assign w1830 = w483 & w1582;
assign w1831 = w483 | w1582;
assign w1832 = w1322 ~^ w1586;
assign w1833 = w1322 ~| w1586;
assign w1834 = w1322 & w1586;
assign w1835 = w1559 ~| w1587;
assign w1836 = w1572 ~^ w1588;
assign w1837 = w1572 | w1588;
assign w1838 = w1572 & w1588;
assign w1839 = w901 ^ w1589;
assign w1840 = w902 ~| w1589;
assign w1841 = w1308 ~^ w1591;
assign w1842 = w1308 ~| w1591;
assign w1843 = ~w1591;
assign w1844 = w898 ~^ w1592;
assign w1845 = w900 | w1592;
assign w1846 = w1584 ~^ w1593;
assign w1847 = w1584 ~| w1595;
assign w1848 = w1585 ~^ w1596;
assign w1849 = w1585 & w1596;
assign w1850 = w1585 | w1596;
assign w1851 = w1368 ~^ w1597;
assign w1852 = ~w1597;
assign w1853 = w960 | w1598;
assign w1854 = w499 | w1600;
assign w1855 = w536 | w1601;
assign w1856 = w1354 ~^ w1602;
assign w1857 = w926 & w1603;
assign w1858 = w926 ~| w1603;
assign w1859 = w923 | w1606;
assign w1860 = w72 & w1609;
assign w1861 = w1604 ~^ w1611;
assign w1862 = w1605 | w1611;
assign w1863 = w931 ~^ w1613;
assign w1864 = w931 | w1613;
assign w1865 = w931 & w1613;
assign w1866 = w1352 ~^ w1614;
assign w1867 = w1352 ~| w1614;
assign w1868 = ~w1614;
assign w1869 = w1349 ~^ w1615;
assign w1870 = w507 ~^ w1616;
assign w1871 = w932 | w1616;
assign w1872 = ~w1616;
assign w1873 = w553 ~^ w1617;
assign w1874 = w553 & w1617;
assign w1875 = w553 | w1617;
assign w1876 = w1362 ~^ w1621;
assign w1877 = w1362 ~| w1621;
assign w1878 = w1362 & w1621;
assign w1879 = w1597 ~| w1622;
assign w1880 = w1607 ~^ w1623;
assign w1881 = w1607 | w1623;
assign w1882 = w1607 & w1623;
assign w1883 = w975 ^ w1624;
assign w1884 = w976 ~| w1624;
assign w1885 = w1348 ~^ w1626;
assign w1886 = w1348 ~| w1626;
assign w1887 = ~w1626;
assign w1888 = w972 ~^ w1627;
assign w1889 = w974 | w1627;
assign w1890 = w1619 ~^ w1628;
assign w1891 = w1619 ~| w1630;
assign w1892 = w1620 ~^ w1631;
assign w1893 = w1620 & w1631;
assign w1894 = w1620 | w1631;
assign w1895 = w1464 & w1633;
assign w1896 = w1464 ~| w1633;
assign w1897 = w1379 | w1634;
assign w1898 = w1413 ~^ w1635;
assign w1899 = ~w1635;
assign w1900 = w1034 | w1636;
assign w1901 = w569 | w1638;
assign w1902 = w606 | w1639;
assign w1903 = w1398 ~^ w1640;
assign w1904 = w1000 & w1641;
assign w1905 = w1000 ~| w1641;
assign w1906 = w997 | w1644;
assign w1907 = w1521 ~^ w1645;
assign w1908 = w1521 & w1646;
assign w1909 = w142 & w1650;
assign w1910 = w1642 ~^ w1652;
assign w1911 = w1643 | w1652;
assign w1912 = w1005 ~^ w1654;
assign w1913 = w1005 | w1654;
assign w1914 = w1005 & w1654;
assign w1915 = w1396 ~^ w1655;
assign w1916 = w1396 ~| w1655;
assign w1917 = ~w1655;
assign w1918 = w1393 ~^ w1656;
assign w1919 = w577 ~^ w1657;
assign w1920 = w1006 | w1657;
assign w1921 = ~w1657;
assign w1922 = w623 ~^ w1658;
assign w1923 = w623 & w1658;
assign w1924 = w623 | w1658;
assign w1925 = w1406 ~^ w1662;
assign w1926 = w1406 ~| w1662;
assign w1927 = w1406 & w1662;
assign w1928 = w1635 ~| w1663;
assign w1929 = w1648 ~^ w1664;
assign w1930 = w1648 | w1664;
assign w1931 = w1648 & w1664;
assign w1932 = w1050 ^ w1665;
assign w1933 = w1051 ~| w1665;
assign w1934 = w1392 ~^ w1667;
assign w1935 = w1392 ~| w1667;
assign w1936 = ~w1667;
assign w1937 = w1047 ~^ w1668;
assign w1938 = w1049 | w1668;
assign w1939 = w1660 ~^ w1669;
assign w1940 = w1660 ~| w1671;
assign w1941 = w1661 ~^ w1672;
assign w1942 = w1661 & w1672;
assign w1943 = w1661 | w1672;
assign w1944 = w1558 & w1674;
assign w1945 = w1456 ~^ w1675;
assign w1946 = ~w1675;
assign w1947 = w1109 | w1676;
assign w1948 = w639 | w1678;
assign w1949 = w676 | w1679;
assign w1950 = ~w1680;
assign w1951 = w1442 ~^ w1681;
assign w1952 = w1075 & w1682;
assign w1953 = w1075 ~| w1682;
assign w1954 = w1072 | w1685;
assign w1955 = w1151 ^ w1686;
assign w1956 = w1151 & w1688;
assign w1957 = w352 | w1690;
assign w1958 = w1649 ~^ w1692;
assign w1959 = w1649 & w1692;
assign w1960 = w1649 | w1692;
assign w1961 = w227 & w1693;
assign w1962 = w1683 ~^ w1695;
assign w1963 = w1684 | w1695;
assign w1964 = w1080 ~^ w1697;
assign w1965 = w1080 | w1697;
assign w1966 = w1080 & w1697;
assign w1967 = w1440 ~^ w1698;
assign w1968 = w1440 ~| w1698;
assign w1969 = ~w1698;
assign w1970 = w1437 ~^ w1699;
assign w1971 = w647 ~^ w1700;
assign w1972 = w1081 | w1700;
assign w1973 = ~w1700;
assign w1974 = w693 ~^ w1701;
assign w1975 = w693 & w1701;
assign w1976 = w693 | w1701;
assign w1977 = w1450 ~^ w1705;
assign w1978 = w1450 ~| w1705;
assign w1979 = w1450 & w1705;
assign w1980 = w1675 ~| w1706;
assign w1981 = w1691 ~^ w1707;
assign w1982 = w1691 | w1707;
assign w1983 = w1691 & w1707;
assign w1984 = w1125 ^ w1708;
assign w1985 = w1126 ~| w1708;
assign w1986 = w1436 ~^ w1710;
assign w1987 = w1436 ~| w1710;
assign w1988 = ~w1710;
assign w1989 = w1122 ~^ w1711;
assign w1990 = w1124 | w1711;
assign w1991 = w1703 ~^ w1712;
assign w1992 = w1703 ~| w1714;
assign w1993 = w1704 ~^ w1715;
assign w1994 = w1704 & w1715;
assign w1995 = w1704 | w1715;
assign w1996 = w1497 ~^ w1717;
assign w1997 = ~w1717;
assign w1998 = w1184 | w1718;
assign w1999 = w709 | w1720;
assign w2000 = w746 | w1721;
assign w2001 = w1483 ~^ w1722;
assign w2002 = w1150 & w1723;
assign w2003 = w1150 ~| w1723;
assign w2004 = w1147 | w1726;
assign w2005 = w1001 ~^ w1727;
assign w2006 = w1001 & w1728;
assign w2007 = w1608 ^ w1730;
assign w2008 = w1608 & w1731;
assign w2009 = w336 & w1735;
assign w2010 = w1724 ~^ w1737;
assign w2011 = w1725 | w1737;
assign w2012 = w1155 ~^ w1739;
assign w2013 = w1155 | w1739;
assign w2014 = w1155 & w1739;
assign w2015 = w1481 ~^ w1740;
assign w2016 = w1481 ~| w1740;
assign w2017 = ~w1740;
assign w2018 = w1478 ~^ w1741;
assign w2019 = w717 ~^ w1742;
assign w2020 = w1156 | w1742;
assign w2021 = ~w1742;
assign w2022 = w763 ~^ w1743;
assign w2023 = w763 & w1743;
assign w2024 = w763 | w1743;
assign w2025 = w1491 ~^ w1747;
assign w2026 = w1491 ~| w1747;
assign w2027 = w1491 & w1747;
assign w2028 = w1717 ~| w1748;
assign w2029 = w1733 ~^ w1749;
assign w2030 = w1733 | w1749;
assign w2031 = w1733 & w1749;
assign w2032 = w1199 ^ w1750;
assign w2033 = w1200 ~| w1750;
assign w2034 = w1477 ~^ w1752;
assign w2035 = w1477 ~| w1752;
assign w2036 = ~w1752;
assign w2037 = w1196 ~^ w1753;
assign w2038 = w1198 | w1753;
assign w2039 = w1745 ~^ w1754;
assign w2040 = w1745 ~| w1756;
assign w2041 = w1746 ~^ w1757;
assign w2042 = w1746 & w1757;
assign w2043 = w1746 | w1757;
assign w2044 = w1555 ~^ w1759;
assign w2045 = w1716 & w1759;
assign w2046 = w1716 | w1759;
assign w2047 = w1632 & w1760;
assign w2048 = w1673 ^ w1761;
assign w2049 = w1511 | w1762;
assign w2050 = w1761 & w1763;
assign w2051 = w1761 ~| w1763;
assign w2052 = w1513 | w1764;
assign w2053 = w1547 ~^ w1765;
assign w2054 = ~w1765;
assign w2055 = w1260 | w1766;
assign w2056 = w779 | w1768;
assign w2057 = w816 | w1769;
assign w2058 = w1532 ~^ w1770;
assign w2059 = w1226 & w1771;
assign w2060 = w1226 ~| w1771;
assign w2061 = w1223 | w1774;
assign w2062 = w1344 ~^ w1775;
assign w2063 = w1344 & w1777;
assign w2064 = w1573 ~^ w1779;
assign w2065 = w1573 ~| w1779;
assign w2066 = ~w1779;
assign w2067 = w355 & w1780;
assign w2068 = w1772 ~^ w1782;
assign w2069 = w1773 | w1782;
assign w2070 = w1231 ~^ w1784;
assign w2071 = w1231 | w1784;
assign w2072 = w1231 & w1784;
assign w2073 = w1530 ~^ w1785;
assign w2074 = w1530 ~| w1785;
assign w2075 = ~w1785;
assign w2076 = w1527 ~^ w1786;
assign w2077 = w787 ~^ w1787;
assign w2078 = w1232 | w1787;
assign w2079 = ~w1787;
assign w2080 = w833 ~^ w1788;
assign w2081 = w833 & w1788;
assign w2082 = w833 | w1788;
assign w2083 = w1540 ~^ w1793;
assign w2084 = w1540 ~| w1793;
assign w2085 = w1540 & w1793;
assign w2086 = w1765 ~| w1794;
assign w2087 = w1778 ~^ w1795;
assign w2088 = w1778 | w1795;
assign w2089 = w1778 & w1795;
assign w2090 = w1277 ^ w1796;
assign w2091 = w1278 ~| w1796;
assign w2092 = w1526 ~^ w1798;
assign w2093 = w1526 ~| w1798;
assign w2094 = ~w1798;
assign w2095 = w1274 ~^ w1799;
assign w2096 = w1276 | w1799;
assign w2097 = w1790 ~^ w1800;
assign w2098 = w1790 ~| w1802;
assign w2099 = w1791 ~^ w1803;
assign w2100 = w1791 & w1803;
assign w2101 = w1791 | w1803;
assign w2102 = w1328 | w1805;
assign w2103 = w1331 ~^ w1806;
assign w2104 = w1590 ~| w1806;
assign w2105 = ~w1806;
assign w2106 = w1807 & w1808;
assign w2107 = w10 & w1809;
assign w2108 = w1314 ~| w1810;
assign w2109 = w1570 | w1814;
assign w2110 = in5[4] & w1816;
assign w2111 = in5[4] | w1816;
assign w2112 = ~w1817;
assign w2113 = w1812 & w1818;
assign w2114 = w1310 ~^ w1819;
assign w2115 = w1310 | w1821;
assign w2116 = w1561 ~^ w1822;
assign w2117 = w1577 | w1824;
assign w2118 = w1323 ~^ w1826;
assign w2119 = w437 ~| w1828;
assign w2120 = w1320 ~^ w1829;
assign w2121 = w1320 | w1830;
assign w2122 = w1317 ~^ w1836;
assign w2123 = w1317 | w1838;
assign w2124 = w2 & w1839;
assign w2125 = w903 | w1840;
assign w2126 = w1575 | w1843;
assign w2127 = w1825 ~^ w1844;
assign w2128 = w1309 | w1844;
assign w2129 = w1309 & w1844;
assign w2130 = w899 & w1845;
assign w2131 = w1594 | w1847;
assign w2132 = w1297 ~^ w1848;
assign w2133 = w1297 | w1849;
assign w2134 = w1368 | w1852;
assign w2135 = w1371 ~^ w1853;
assign w2136 = w1625 ~| w1853;
assign w2137 = ~w1853;
assign w2138 = w1854 & w1855;
assign w2139 = w80 & w1856;
assign w2140 = w1354 ~| w1857;
assign w2141 = ~w1860;
assign w2142 = ~w1861;
assign w2143 = w1859 & w1862;
assign w2144 = w1350 ~^ w1863;
assign w2145 = w1350 | w1865;
assign w2146 = w1599 ~^ w1866;
assign w2147 = w1612 | w1868;
assign w2148 = w1363 ~^ w1870;
assign w2149 = w507 ~| w1872;
assign w2150 = w1360 ~^ w1873;
assign w2151 = w1360 | w1874;
assign w2152 = w1357 ~^ w1880;
assign w2153 = w1357 | w1882;
assign w2154 = w72 & w1883;
assign w2155 = w977 | w1884;
assign w2156 = w1610 | w1887;
assign w2157 = w1869 ~^ w1888;
assign w2158 = w1349 | w1888;
assign w2159 = w1349 & w1888;
assign w2160 = w973 & w1889;
assign w2161 = w1629 | w1891;
assign w2162 = w1337 ~^ w1892;
assign w2163 = w1337 | w1893;
assign w2164 = w1413 | w1899;
assign w2165 = w1416 ~^ w1900;
assign w2166 = w1666 ~| w1900;
assign w2167 = ~w1900;
assign w2168 = w1901 & w1902;
assign w2169 = w150 & w1903;
assign w2170 = w1398 ~| w1904;
assign w2171 = w1897 ~| w1907;
assign w2172 = w1897 & w1907;
assign w2173 = w1647 | w1908;
assign w2174 = ~w1910;
assign w2175 = w1906 & w1911;
assign w2176 = w1394 ~^ w1912;
assign w2177 = w1394 | w1914;
assign w2178 = w1637 ~^ w1915;
assign w2179 = w1653 | w1917;
assign w2180 = w1407 ~^ w1919;
assign w2181 = w577 ~| w1921;
assign w2182 = w1404 ~^ w1922;
assign w2183 = w1404 | w1923;
assign w2184 = w1401 ~^ w1929;
assign w2185 = w1401 | w1931;
assign w2186 = w142 & w1932;
assign w2187 = w1052 | w1933;
assign w2188 = w1651 | w1936;
assign w2189 = w1918 ~^ w1937;
assign w2190 = w1393 | w1937;
assign w2191 = w1393 & w1937;
assign w2192 = w1048 & w1938;
assign w2193 = w1670 | w1940;
assign w2194 = w1381 ~^ w1941;
assign w2195 = w1381 | w1942;
assign w2196 = w1456 | w1946;
assign w2197 = w1459 ~^ w1947;
assign w2198 = w1709 ~| w1947;
assign w2199 = ~w1947;
assign w2200 = w1948 & w1949;
assign w2201 = w235 & w1951;
assign w2202 = w1442 ~| w1952;
assign w2203 = w1897 ^ w1955;
assign w2204 = w1687 | w1956;
assign w2205 = w1860 ~^ w1957;
assign w2206 = ~w1957;
assign w2207 = w1734 ~^ w1958;
assign w2208 = w1734 & w1960;
assign w2209 = w1961 ~^ in5[4];
assign w2210 = ~w1962;
assign w2211 = w1954 & w1963;
assign w2212 = w1438 ~^ w1964;
assign w2213 = w1438 | w1966;
assign w2214 = w1677 ~^ w1967;
assign w2215 = w1696 | w1969;
assign w2216 = w1451 ~^ w1971;
assign w2217 = w647 ~| w1973;
assign w2218 = w1448 ~^ w1974;
assign w2219 = w1448 | w1975;
assign w2220 = w1445 ~^ w1981;
assign w2221 = w1445 | w1983;
assign w2222 = w227 & w1984;
assign w2223 = w1127 | w1985;
assign w2224 = w1694 | w1988;
assign w2225 = w1970 ~^ w1989;
assign w2226 = w1437 | w1989;
assign w2227 = w1437 & w1989;
assign w2228 = w1123 & w1990;
assign w2229 = w1713 | w1992;
assign w2230 = w1423 ~^ w1993;
assign w2231 = w1423 | w1994;
assign w2232 = w1497 | w1997;
assign w2233 = w1500 ~^ w1998;
assign w2234 = w1751 ~| w1998;
assign w2235 = ~w1998;
assign w2236 = w1999 & w2000;
assign w2237 = w344 & w2001;
assign w2238 = w1483 ~| w2002;
assign w2239 = w1813 ~^ w2005;
assign w2240 = ~w2005;
assign w2241 = w1729 | w2006;
assign w2242 = w1732 | w2008;
assign w2243 = w1909 ~^ w2009;
assign w2244 = ~w2010;
assign w2245 = w2004 & w2011;
assign w2246 = w1479 ~^ w2012;
assign w2247 = w1479 | w2014;
assign w2248 = w1719 ~^ w2015;
assign w2249 = w1738 | w2017;
assign w2250 = w1492 ~^ w2019;
assign w2251 = w717 ~| w2021;
assign w2252 = w1489 ~^ w2022;
assign w2253 = w1489 | w2023;
assign w2254 = w1486 ~^ w2029;
assign w2255 = w1486 | w2031;
assign w2256 = w336 & w2032;
assign w2257 = w1201 | w2033;
assign w2258 = w1736 | w2036;
assign w2259 = w2018 ~^ w2037;
assign w2260 = w1478 | w2037;
assign w2261 = w1478 & w2037;
assign w2262 = w1197 & w2038;
assign w2263 = w1755 | w2040;
assign w2264 = w1466 ~^ w2041;
assign w2265 = w1466 | w2042;
assign out1[0] = w1716 ~^ w2044;
assign w2266 = w1555 & w2046;
assign w2267 = w1896 ~| w2047;
assign w2268 = w1464 ^ w2047;
assign w2269 = w1763 ~^ w2048;
assign w2270 = w1944 ^ w2049;
assign w2271 = w1673 ~| w2051;
assign w2272 = w2049 & w2052;
assign w2273 = w2049 ~| w2052;
assign w2274 = w1547 | w2054;
assign w2275 = w1550 ~^ w2055;
assign w2276 = w1797 ~| w2055;
assign w2277 = ~w2055;
assign w2278 = w2056 & w2057;
assign w2279 = w363 & w2058;
assign w2280 = w1532 ~| w2059;
assign w2281 = w1776 | w2063;
assign w2282 = w1689 ~^ w2064;
assign w2283 = w1689 | w2065;
assign w2284 = w1815 | w2066;
assign w2285 = w2009 | w2067;
assign w2286 = w2009 & w2067;
assign w2287 = ~w2068;
assign w2288 = w2061 & w2069;
assign w2289 = w1528 ~^ w2070;
assign w2290 = w1528 | w2072;
assign w2291 = w1767 ~^ w2073;
assign w2292 = w1783 | w2075;
assign w2293 = w1541 ~^ w2077;
assign w2294 = w787 ~| w2079;
assign w2295 = w1538 ~^ w2080;
assign w2296 = w1538 | w2081;
assign w2297 = w1535 ~^ w2087;
assign w2298 = w1535 | w2089;
assign w2299 = w355 & w2090;
assign w2300 = w1279 | w2091;
assign w2301 = w1781 | w2094;
assign w2302 = w2076 ~^ w2095;
assign w2303 = w1527 | w2095;
assign w2304 = w1527 & w2095;
assign w2305 = w1275 & w2096;
assign w2306 = w1801 | w2098;
assign w2307 = w1515 ~^ w2099;
assign w2308 = w1515 | w2100;
assign w2309 = w1331 | w2105;
assign w2310 = w1324 ~^ w2106;
assign w2311 = w1583 ~| w2106;
assign w2312 = w1583 & w2106;
assign w2313 = w1811 | w2108;
assign w2314 = ~w2109;
assign w2315 = w1961 & w2111;
assign w2316 = w1804 ~^ w2113;
assign w2317 = w1835 | w2113;
assign w2318 = w1820 & w2115;
assign w2319 = w11 & w2116;
assign w2320 = w1561 & w2117;
assign w2321 = w1841 ~^ w2118;
assign w2322 = w1323 | w2119;
assign w2323 = w1831 & w2121;
assign w2324 = ~w2122;
assign w2325 = w1837 & w2123;
assign w2326 = w13 & w2125;
assign w2327 = w2118 & w2126;
assign w2328 = ~w2127;
assign w2329 = w1580 | w2129;
assign w2330 = w2120 ~^ w2130;
assign w2331 = w2120 ~| w2130;
assign w2332 = w2120 & w2130;
assign w2333 = ~w2131;
assign w2334 = ~w2132;
assign w2335 = w1850 & w2133;
assign w2336 = w1371 | w2137;
assign w2337 = w1364 ~^ w2138;
assign w2338 = w1618 ~| w2138;
assign w2339 = w1618 & w2138;
assign w2340 = ~w2139;
assign w2341 = w1858 | w2140;
assign w2342 = w1957 ~| w2141;
assign w2343 = w1851 ~^ w2143;
assign w2344 = w1879 | w2143;
assign w2345 = w1864 & w2145;
assign w2346 = w81 & w2146;
assign w2347 = w1599 & w2147;
assign w2348 = w1885 ~^ w2148;
assign w2349 = w1363 | w2149;
assign w2350 = w1875 & w2151;
assign w2351 = ~w2152;
assign w2352 = w1881 & w2153;
assign w2353 = w83 & w2155;
assign w2354 = w2148 & w2156;
assign w2355 = ~w2157;
assign w2356 = w1615 | w2159;
assign w2357 = w2150 ~^ w2160;
assign w2358 = w2150 ~| w2160;
assign w2359 = w2150 & w2160;
assign w2360 = ~w2161;
assign w2361 = ~w2162;
assign w2362 = w1894 & w2163;
assign w2363 = w1416 | w2167;
assign w2364 = w1408 ~^ w2168;
assign w2365 = w1659 ~| w2168;
assign w2366 = w1659 & w2168;
assign w2367 = w2139 ~| w2169;
assign w2368 = ~w2169;
assign w2369 = w1905 | w2170;
assign w2370 = w1955 ~| w2171;
assign w2371 = w1680 ~^ w2173;
assign w2372 = w1898 ~^ w2175;
assign w2373 = w1928 | w2175;
assign w2374 = w1913 & w2177;
assign w2375 = w151 & w2178;
assign w2376 = w1637 & w2179;
assign w2377 = w1934 ~^ w2180;
assign w2378 = w1407 | w2181;
assign w2379 = w1924 & w2183;
assign w2380 = ~w2184;
assign w2381 = w1930 & w2185;
assign w2382 = w2154 ~^ w2186;
assign w2383 = w2154 & w2186;
assign w2384 = w2154 | w2186;
assign w2385 = w153 & w2187;
assign w2386 = w2180 & w2188;
assign w2387 = ~w2189;
assign w2388 = w1656 | w2191;
assign w2389 = w2182 ~^ w2192;
assign w2390 = w2182 ~| w2192;
assign w2391 = w2182 & w2192;
assign w2392 = ~w2193;
assign w2393 = ~w2194;
assign w2394 = w1943 & w2195;
assign w2395 = w1459 | w2199;
assign w2396 = w1452 ~^ w2200;
assign w2397 = w1702 ~| w2200;
assign w2398 = w1702 & w2200;
assign w2399 = w1953 | w2202;
assign w2400 = w1907 ~^ w2203;
assign w2401 = w1950 | w2204;
assign w2402 = ~w2204;
assign w2403 = w1860 | w2206;
assign w2404 = w2109 ~^ w2207;
assign w2405 = ~w2207;
assign w2406 = w1959 | w2208;
assign w2407 = w1816 ~^ w2209;
assign w2408 = w1945 ~^ w2211;
assign w2409 = w1980 | w2211;
assign w2410 = w1965 & w2213;
assign w2411 = w236 & w2214;
assign w2412 = w1677 & w2215;
assign w2413 = w1986 ~^ w2216;
assign w2414 = w1451 | w2217;
assign w2415 = w1976 & w2219;
assign w2416 = ~w2220;
assign w2417 = w1982 & w2221;
assign w2418 = ~w2222;
assign w2419 = w238 & w2223;
assign w2420 = w2216 & w2224;
assign w2421 = ~w2225;
assign w2422 = w1699 | w2227;
assign w2423 = w2218 ~^ w2228;
assign w2424 = w2218 ~| w2228;
assign w2425 = w2218 & w2228;
assign w2426 = ~w2229;
assign w2427 = ~w2230;
assign w2428 = w1995 & w2231;
assign w2429 = w1500 | w2235;
assign w2430 = w1493 ~^ w2236;
assign w2431 = w1744 ~| w2236;
assign w2432 = w1744 & w2236;
assign w2433 = w2201 ~^ w2237;
assign w2434 = w2107 & w2237;
assign w2435 = w2107 | w2237;
assign w2436 = w2003 | w2238;
assign w2437 = ~w2239;
assign w2438 = w1813 | w2240;
assign w2439 = w2007 ^ w2241;
assign w2440 = w2062 ~| w2241;
assign w2441 = w2062 & w2241;
assign w2442 = w2067 ~^ w2243;
assign w2443 = w1996 ~^ w2245;
assign w2444 = w2028 | w2245;
assign w2445 = w2013 & w2247;
assign w2446 = w345 & w2248;
assign w2447 = w1719 & w2249;
assign w2448 = w2034 ~^ w2250;
assign w2449 = w1492 | w2251;
assign w2450 = w2024 & w2253;
assign w2451 = ~w2254;
assign w2452 = w2030 & w2255;
assign w2453 = w2222 ~^ w2256;
assign w2454 = ~w2256;
assign w2455 = w347 & w2257;
assign w2456 = w2250 & w2258;
assign w2457 = ~w2259;
assign w2458 = w1741 | w2261;
assign w2459 = w2252 ~^ w2262;
assign w2460 = w2252 ~| w2262;
assign w2461 = w2252 & w2262;
assign w2462 = ~w2263;
assign w2463 = ~w2264;
assign w2464 = w2043 & w2265;
assign w2465 = w2045 | w2266;
assign w2466 = w1895 | w2267;
assign w2467 = w1633 ~^ w2268;
assign w2468 = w2052 ~^ w2270;
assign w2469 = w2050 | w2271;
assign w2470 = w1944 ~| w2273;
assign w2471 = w1550 | w2277;
assign w2472 = w1542 ~^ w2278;
assign w2473 = w1789 ~| w2278;
assign w2474 = w1789 & w2278;
assign w2475 = w2169 ~^ w2279;
assign w2476 = ~w2279;
assign w2477 = w2060 | w2280;
assign w2478 = w2205 ~^ w2281;
assign w2479 = w2283 & w2284;
assign w2480 = w1909 & w2285;
assign w2481 = w2053 ~^ w2288;
assign w2482 = w2086 | w2288;
assign w2483 = w2071 & w2290;
assign w2484 = w364 & w2291;
assign w2485 = w1767 & w2292;
assign w2486 = w2092 ~^ w2293;
assign w2487 = w1541 | w2294;
assign w2488 = w2082 & w2296;
assign w2489 = ~w2297;
assign w2490 = w2088 & w2298;
assign w2491 = w366 & w2300;
assign w2492 = w2293 & w2301;
assign w2493 = ~w2302;
assign w2494 = w1786 | w2304;
assign w2495 = w2295 ~^ w2305;
assign w2496 = w2295 ~| w2305;
assign w2497 = w2295 & w2305;
assign w2498 = ~w2306;
assign w2499 = ~w2307;
assign w2500 = w2101 & w2308;
assign w2501 = w2114 ~^ w2310;
assign w2502 = w2114 ~| w2312;
assign w2503 = w3 & w2313;
assign w2504 = w2110 | w2315;
assign w2505 = w2102 & w2317;
assign w2506 = w1817 ~^ w2318;
assign w2507 = w2112 & w2318;
assign w2508 = w2112 ~| w2318;
assign w2509 = w1823 | w2320;
assign w2510 = ~w2321;
assign w2511 = w1827 & w2322;
assign w2512 = w1832 ^ w2323;
assign w2513 = w1834 ~| w2323;
assign w2514 = ~w2324;
assign w2515 = w2321 ~^ w2325;
assign w2516 = w1842 | w2327;
assign w2517 = w2128 & w2329;
assign w2518 = w2132 ~^ w2333;
assign w2519 = w2132 ~| w2333;
assign w2520 = w2131 | w2334;
assign w2521 = w2103 ~^ w2335;
assign w2522 = w2104 | w2335;
assign w2523 = w2144 ~^ w2337;
assign w2524 = w2144 ~| w2339;
assign w2525 = w73 & w2341;
assign w2526 = w2134 & w2344;
assign w2527 = w1861 ~^ w2345;
assign w2528 = w2142 & w2345;
assign w2529 = w2142 ~| w2345;
assign w2530 = w1867 | w2347;
assign w2531 = ~w2348;
assign w2532 = w1871 & w2349;
assign w2533 = w1876 ^ w2350;
assign w2534 = w1878 ~| w2350;
assign w2535 = ~w2351;
assign w2536 = w2348 ~^ w2352;
assign w2537 = w1505 ~^ w2353;
assign w2538 = w484 & w2353;
assign w2539 = w484 ~| w2353;
assign w2540 = w1886 | w2354;
assign w2541 = w2158 & w2356;
assign w2542 = w2162 ~^ w2360;
assign w2543 = w2162 ~| w2360;
assign w2544 = w2161 | w2361;
assign w2545 = w2135 ~^ w2362;
assign w2546 = w2136 | w2362;
assign w2547 = w2176 ~^ w2364;
assign w2548 = w2176 ~| w2366;
assign w2549 = w2340 | w2368;
assign w2550 = w143 & w2369;
assign w2551 = w2172 | w2370;
assign w2552 = w2204 ~^ w2371;
assign w2553 = w2164 & w2373;
assign w2554 = w1910 ~^ w2374;
assign w2555 = w2174 & w2374;
assign w2556 = w2174 ~| w2374;
assign w2557 = w1916 | w2376;
assign w2558 = ~w2377;
assign w2559 = w1920 & w2378;
assign w2560 = w1925 ^ w2379;
assign w2561 = w1927 ~| w2379;
assign w2562 = ~w2380;
assign w2563 = w2377 ~^ w2381;
assign w2564 = w2299 ~^ w2382;
assign w2565 = w2299 & w2384;
assign w2566 = w2326 ~^ w2385;
assign w2567 = w1935 | w2386;
assign w2568 = w2190 & w2388;
assign w2569 = w2194 ~^ w2392;
assign w2570 = w2194 ~| w2392;
assign w2571 = w2193 | w2393;
assign w2572 = w2165 ~^ w2394;
assign w2573 = w2166 | w2394;
assign w2574 = w2212 ~^ w2396;
assign w2575 = w2212 ~| w2398;
assign w2576 = w228 & w2399;
assign w2577 = ~w2400;
assign w2578 = w2173 & w2401;
assign w2579 = w1680 ~| w2402;
assign w2580 = w2281 & w2403;
assign w2581 = w2282 ~^ w2404;
assign w2582 = w2282 | w2405;
assign w2583 = w2282 & w2405;
assign w2584 = w2242 ~^ w2406;
assign w2585 = w2242 & w2406;
assign w2586 = w2242 | w2406;
assign w2587 = ~w2407;
assign w2588 = w2196 & w2409;
assign w2589 = w1962 ~^ w2410;
assign w2590 = w2210 & w2410;
assign w2591 = w2210 ~| w2410;
assign w2592 = w2319 | w2411;
assign w2593 = w2319 & w2411;
assign w2594 = w1968 | w2412;
assign w2595 = ~w2413;
assign w2596 = w1972 & w2414;
assign w2597 = w1977 ^ w2415;
assign w2598 = w1979 ~| w2415;
assign w2599 = ~w2416;
assign w2600 = w2413 ~^ w2417;
assign w2601 = w2385 | w2419;
assign w2602 = w2385 & w2419;
assign w2603 = w1987 | w2420;
assign w2604 = w2226 & w2422;
assign w2605 = w2230 ~^ w2426;
assign w2606 = w2230 ~| w2426;
assign w2607 = w2229 | w2427;
assign w2608 = w2197 ~^ w2428;
assign w2609 = w2198 | w2428;
assign w2610 = w2246 ~^ w2430;
assign w2611 = w2246 ~| w2432;
assign w2612 = w2107 ~^ w2433;
assign w2613 = w2201 & w2435;
assign w2614 = w337 & w2436;
assign w2615 = w2400 ~^ w2437;
assign w2616 = ~w2437;
assign w2617 = w2062 ~^ w2439;
assign w2618 = w2007 ~| w2440;
assign w2619 = ~w2442;
assign w2620 = w2232 & w2444;
assign w2621 = w2010 ~^ w2445;
assign w2622 = w2244 & w2445;
assign w2623 = w2244 ~| w2445;
assign w2624 = w2411 ~^ w2446;
assign w2625 = w2016 | w2447;
assign w2626 = ~w2448;
assign w2627 = w2020 & w2449;
assign w2628 = w2025 ^ w2450;
assign w2629 = w2027 ~| w2450;
assign w2630 = ~w2451;
assign w2631 = w2448 ~^ w2452;
assign w2632 = w2124 ~^ w2453;
assign w2633 = w2418 | w2454;
assign w2634 = w2035 | w2456;
assign w2635 = w2260 & w2458;
assign w2636 = w2264 ~^ w2462;
assign w2637 = w2264 ~| w2462;
assign w2638 = w2263 | w2463;
assign w2639 = w2233 ~^ w2464;
assign w2640 = w2234 | w2464;
assign w2641 = w1556 ~^ w2467;
assign w2642 = w1070 ~| w2467;
assign w2643 = w1070 & w2467;
assign w2644 = w2468 ~^ w2469;
assign w2645 = w2468 & w2469;
assign w2646 = w2468 | w2469;
assign w2647 = w2272 | w2470;
assign w2648 = w2289 ~^ w2472;
assign w2649 = w2289 ~| w2474;
assign w2650 = w2139 ~^ w2475;
assign w2651 = w2367 | w2476;
assign w2652 = w356 & w2477;
assign w2653 = ~w2478;
assign w2654 = w2407 ~^ w2479;
assign w2655 = w2286 | w2480;
assign w2656 = w2274 & w2482;
assign w2657 = w2068 ~^ w2483;
assign w2658 = w2287 & w2483;
assign w2659 = w2287 ~| w2483;
assign w2660 = w2074 | w2485;
assign w2661 = ~w2486;
assign w2662 = w2078 & w2487;
assign w2663 = w2083 ^ w2488;
assign w2664 = w2085 ~| w2488;
assign w2665 = ~w2489;
assign w2666 = w2486 ~^ w2490;
assign w2667 = w2455 ~^ w2491;
assign w2668 = w2455 & w2491;
assign w2669 = w2455 ~| w2491;
assign w2670 = w2093 | w2492;
assign w2671 = w2303 & w2494;
assign w2672 = w2307 ~^ w2498;
assign w2673 = w2307 ~| w2498;
assign w2674 = w2306 | w2499;
assign w2675 = w2275 ~^ w2500;
assign w2676 = w2276 | w2500;
assign w2677 = w11 & w2501;
assign w2678 = w2311 | w2502;
assign w2679 = w2122 ~^ w2505;
assign w2680 = ~w2505;
assign w2681 = w1846 ~^ w2506;
assign w2682 = w1846 ~| w2507;
assign w2683 = w3 & w2509;
assign w2684 = w2325 ~| w2510;
assign w2685 = w2325 & w2510;
assign w2686 = w2127 ~^ w2511;
assign w2687 = w2127 ~| w2511;
assign w2688 = ~w2511;
assign w2689 = w4 & w2512;
assign w2690 = w1833 | w2513;
assign w2691 = w2505 ~| w2514;
assign w2692 = w2330 ^ w2517;
assign w2693 = w2332 ~| w2517;
assign w2694 = w2316 ~^ w2518;
assign w2695 = w2316 & w2520;
assign w2696 = w2309 & w2522;
assign w2697 = w81 & w2523;
assign w2698 = w2338 | w2524;
assign w2699 = w2503 ~^ w2525;
assign w2700 = w2152 ~^ w2526;
assign w2701 = ~w2526;
assign w2702 = w1890 ~^ w2527;
assign w2703 = w1890 ~| w2528;
assign w2704 = w73 & w2530;
assign w2705 = w2352 ~| w2531;
assign w2706 = w2352 & w2531;
assign w2707 = w2157 ~^ w2532;
assign w2708 = w2157 ~| w2532;
assign w2709 = ~w2532;
assign w2710 = w74 & w2533;
assign w2711 = w1877 | w2534;
assign w2712 = w2526 ~| w2535;
assign w2713 = w1215 ~| w2539;
assign w2714 = w2357 ^ w2541;
assign w2715 = w2359 ~| w2541;
assign w2716 = w2343 ~^ w2542;
assign w2717 = w2343 & w2544;
assign w2718 = w2336 & w2546;
assign w2719 = w151 & w2547;
assign w2720 = w2365 | w2548;
assign w2721 = w2346 ~^ w2550;
assign w2722 = w2375 | w2550;
assign w2723 = w2375 & w2550;
assign w2724 = ~w2551;
assign w2725 = ~w2552;
assign w2726 = w2184 ~^ w2553;
assign w2727 = ~w2553;
assign w2728 = w1939 ~^ w2554;
assign w2729 = w1939 ~| w2555;
assign w2730 = w143 & w2557;
assign w2731 = w2381 ~| w2558;
assign w2732 = w2381 & w2558;
assign w2733 = w2189 ~^ w2559;
assign w2734 = w2189 ~| w2559;
assign w2735 = ~w2559;
assign w2736 = w144 & w2560;
assign w2737 = w1926 | w2561;
assign w2738 = w2553 ~| w2562;
assign w2739 = w2383 | w2565;
assign w2740 = w2419 ~^ w2566;
assign w2741 = w2389 ^ w2568;
assign w2742 = w2391 ~| w2568;
assign w2743 = w2372 ~^ w2569;
assign w2744 = w2372 & w2571;
assign w2745 = w2363 & w2573;
assign w2746 = w236 & w2574;
assign w2747 = w2397 | w2575;
assign w2748 = w2576 ~^ in5[5];
assign w2749 = w2437 ~| w2577;
assign w2750 = w2578 | w2579;
assign w2751 = w2342 | w2580;
assign w2752 = w2314 | w2583;
assign w2753 = ~w2587;
assign w2754 = w2220 ~^ w2588;
assign w2755 = ~w2588;
assign w2756 = w1991 ~^ w2589;
assign w2757 = w1991 ~| w2590;
assign w2758 = w2446 & w2592;
assign w2759 = w228 & w2594;
assign w2760 = w2417 ~| w2595;
assign w2761 = w2417 & w2595;
assign w2762 = w2225 ~^ w2596;
assign w2763 = w2225 ~| w2596;
assign w2764 = ~w2596;
assign w2765 = w229 & w2597;
assign w2766 = w1978 | w2598;
assign w2767 = w2588 ~| w2599;
assign w2768 = w2326 & w2601;
assign w2769 = w2423 ^ w2604;
assign w2770 = w2425 ~| w2604;
assign w2771 = w2408 ~^ w2605;
assign w2772 = w2408 & w2607;
assign w2773 = w2395 & w2609;
assign w2774 = w345 & w2610;
assign w2775 = w2431 | w2611;
assign w2776 = w2584 ~^ w2612;
assign w2777 = w2586 & w2612;
assign w2778 = w2434 | w2613;
assign w2779 = w2503 | w2614;
assign w2780 = w2503 & w2614;
assign w2781 = w2400 | w2616;
assign w2782 = w2438 ^ w2617;
assign w2783 = ~w2617;
assign w2784 = w2441 | w2618;
assign w2785 = w2478 ~| w2619;
assign w2786 = w2254 ~^ w2620;
assign w2787 = ~w2620;
assign w2788 = w2039 ~^ w2621;
assign w2789 = w2039 ~| w2622;
assign w2790 = w2319 ~^ w2624;
assign w2791 = w337 & w2625;
assign w2792 = w2452 ~| w2626;
assign w2793 = w2452 & w2626;
assign w2794 = w2259 ~^ w2627;
assign w2795 = w2259 ~| w2627;
assign w2796 = ~w2627;
assign w2797 = w338 & w2628;
assign w2798 = w2026 | w2629;
assign w2799 = w2620 ~| w2630;
assign w2800 = w2459 ^ w2635;
assign w2801 = w2461 ~| w2635;
assign w2802 = w2443 ~^ w2636;
assign w2803 = w2443 & w2638;
assign w2804 = w2429 & w2640;
assign w2805 = w2269 ~^ w2641;
assign w2806 = w2269 & w2641;
assign w2807 = w2269 | w2641;
assign w2808 = w1557 ~| w2642;
assign w2809 = w2466 ~^ w2644;
assign w2810 = w2466 & w2646;
assign w2811 = w2552 ~^ w2647;
assign w2812 = ~w2647;
assign w2813 = w364 & w2648;
assign w2814 = w2473 | w2649;
assign w2815 = ~w2650;
assign w2816 = w2549 & w2651;
assign w2817 = in5[5] | w2652;
assign w2818 = in5[5] & w2652;
assign w2819 = w2442 | w2653;
assign w2820 = w2650 ~^ w2654;
assign w2821 = ~w2655;
assign w2822 = w2297 ~^ w2656;
assign w2823 = ~w2656;
assign w2824 = w2097 ~^ w2657;
assign w2825 = w2097 ~| w2658;
assign w2826 = w356 & w2660;
assign w2827 = w2490 ~| w2661;
assign w2828 = w2490 & w2661;
assign w2829 = w2302 ~^ w2662;
assign w2830 = w2302 ~| w2662;
assign w2831 = ~w2662;
assign w2832 = w357 & w2663;
assign w2833 = w2084 | w2664;
assign w2834 = w2656 ~| w2665;
assign w2835 = w2633 ~^ w2667;
assign w2836 = w2633 ~| w2669;
assign w2837 = w2495 ^ w2671;
assign w2838 = w2497 ~| w2671;
assign w2839 = w2481 ~^ w2672;
assign w2840 = w2481 & w2674;
assign w2841 = w2471 & w2676;
assign w2842 = w0 & w2678;
assign w2843 = w2521 ~^ w2679;
assign w2844 = w2324 | w2680;
assign w2845 = w8 & w2681;
assign w2846 = w2508 | w2682;
assign w2847 = in5[6] | w2683;
assign w2848 = in5[6] & w2683;
assign w2849 = w2516 ~^ w2686;
assign w2850 = w2328 | w2688;
assign w2851 = w10 & w2690;
assign w2852 = w0 & w2692;
assign w2853 = w2331 | w2693;
assign w2854 = w14 & w2694;
assign w2855 = w2519 | w2695;
assign w2856 = w2515 ~^ w2696;
assign w2857 = w2685 ~| w2696;
assign w2858 = w70 & w2698;
assign w2859 = w2614 ~^ w2699;
assign w2860 = w2545 ~^ w2700;
assign w2861 = w2351 | w2701;
assign w2862 = w78 & w2702;
assign w2863 = w2529 | w2703;
assign w2864 = w2540 ~^ w2707;
assign w2865 = w2355 | w2709;
assign w2866 = w80 & w2711;
assign w2867 = w2538 | w2713;
assign w2868 = w70 & w2714;
assign w2869 = w2358 | w2715;
assign w2870 = w84 & w2716;
assign w2871 = w2543 | w2717;
assign w2872 = w2536 ~^ w2718;
assign w2873 = w2706 ~| w2718;
assign w2874 = w2697 & w2719;
assign w2875 = w2697 | w2719;
assign w2876 = w140 & w2720;
assign w2877 = w2375 ~^ w2721;
assign w2878 = w2346 & w2722;
assign w2879 = w2647 ~| w2725;
assign w2880 = w2572 ~^ w2726;
assign w2881 = w2380 | w2727;
assign w2882 = w148 & w2728;
assign w2883 = w2556 | w2729;
assign w2884 = w2567 ~^ w2733;
assign w2885 = w2387 | w2735;
assign w2886 = w2710 ~^ w2736;
assign w2887 = w2710 | w2736;
assign w2888 = w2710 & w2736;
assign w2889 = w150 & w2737;
assign w2890 = w1411 ~^ w2739;
assign w2891 = w2537 ~^ w2740;
assign w2892 = ~w2740;
assign w2893 = w140 & w2741;
assign w2894 = w2390 | w2742;
assign w2895 = w154 & w2743;
assign w2896 = w2570 | w2744;
assign w2897 = w2563 ~^ w2745;
assign w2898 = w2732 ~| w2745;
assign w2899 = w225 & w2747;
assign w2900 = w2652 ~^ w2748;
assign w2901 = w2442 ~^ w2750;
assign w2902 = w2582 & w2752;
assign w2903 = w2650 ~| w2753;
assign w2904 = w2608 ~^ w2754;
assign w2905 = w2416 | w2755;
assign w2906 = w233 & w2756;
assign w2907 = w2591 | w2757;
assign w2908 = w2593 | w2758;
assign w2909 = w2759 ~^ in5[6];
assign w2910 = w2603 ~^ w2762;
assign w2911 = w2421 | w2764;
assign w2912 = ~w2765;
assign w2913 = w235 & w2766;
assign w2914 = w2602 | w2768;
assign w2915 = w225 & w2769;
assign w2916 = w2424 | w2770;
assign w2917 = w239 & w2771;
assign w2918 = w2606 | w2772;
assign w2919 = w2600 ~^ w2773;
assign w2920 = w2761 ~| w2773;
assign w2921 = w2746 ~^ w2774;
assign w2922 = w2677 & w2774;
assign w2923 = w2677 | w2774;
assign w2924 = w334 & w2775;
assign w2925 = ~w2776;
assign w2926 = w2585 | w2777;
assign w2927 = w2484 ~^ w2778;
assign w2928 = w2484 & w2778;
assign w2929 = w2484 | w2778;
assign w2930 = w2525 & w2779;
assign w2931 = w2581 ~^ w2782;
assign w2932 = w2581 & w2783;
assign w2933 = w2581 ~| w2783;
assign w2934 = w2776 ~| w2784;
assign w2935 = ~w2784;
assign w2936 = w2639 ~^ w2786;
assign w2937 = w2451 | w2787;
assign w2938 = w342 & w2788;
assign w2939 = w2623 | w2789;
assign w2940 = ~w2790;
assign w2941 = w2730 ~^ w2791;
assign w2942 = w2634 ~^ w2794;
assign w2943 = w2457 | w2796;
assign w2944 = w2765 ~^ w2797;
assign w2945 = ~w2797;
assign w2946 = w344 & w2798;
assign w2947 = w334 & w2800;
assign w2948 = w2460 | w2801;
assign w2949 = w348 & w2802;
assign w2950 = w2637 | w2803;
assign w2951 = w2631 ~^ w2804;
assign w2952 = w2793 ~| w2804;
assign out1[1] = w2465 ~^ w2805;
assign w2953 = w2465 & w2807;
assign w2954 = w2643 | w2808;
assign w2955 = ~w2809;
assign w2956 = w2645 | w2810;
assign w2957 = w2551 ~^ w2811;
assign w2958 = w2552 | w2812;
assign w2959 = w2719 ~^ w2813;
assign w2960 = w353 & w2814;
assign w2961 = w2587 | w2815;
assign w2962 = w2576 & w2817;
assign w2963 = w2750 & w2819;
assign w2964 = w2816 ~^ w2821;
assign w2965 = w2675 ~^ w2822;
assign w2966 = w2489 | w2823;
assign w2967 = w361 & w2824;
assign w2968 = w2659 | w2825;
assign w2969 = w2791 & w2826;
assign w2970 = w2791 | w2826;
assign w2971 = w2670 ~^ w2829;
assign w2972 = w2493 | w2831;
assign w2973 = w363 & w2833;
assign w2974 = ~w2835;
assign w2975 = w2668 | w2836;
assign w2976 = w353 & w2837;
assign w2977 = w2496 | w2838;
assign w2978 = w367 & w2839;
assign w2979 = w2673 | w2840;
assign w2980 = w2666 ~^ w2841;
assign w2981 = w2828 ~| w2841;
assign w2982 = w13 & w2843;
assign w2983 = w2521 & w2844;
assign w2984 = w6 & w2846;
assign w2985 = w2759 & w2847;
assign w2986 = w12 & w2849;
assign w2987 = w2516 & w2850;
assign w2988 = w12 & w2853;
assign w2989 = w5 & w2855;
assign w2990 = w9 & w2856;
assign w2991 = w2684 | w2857;
assign w2992 = w2655 ~| w2859;
assign w2993 = ~w2859;
assign w2994 = w83 & w2860;
assign w2995 = w2545 & w2861;
assign w2996 = w2842 ~^ w2862;
assign w2997 = w76 & w2863;
assign w2998 = w82 & w2864;
assign w2999 = w2540 & w2865;
assign w3000 = w2632 ~^ w2866;
assign w3001 = w2124 ~| w2866;
assign w3002 = w2124 & w2866;
assign w3003 = w1792 ~^ w2867;
assign w3004 = w82 & w2869;
assign w3005 = ~w2870;
assign w3006 = w75 & w2871;
assign w3007 = w79 & w2872;
assign w3008 = w2705 | w2873;
assign w3009 = w2813 & w2875;
assign w3010 = w2858 ~^ w2876;
assign w3011 = ~w2877;
assign w3012 = w2723 | w2878;
assign w3013 = w2724 | w2879;
assign w3014 = w153 & w2880;
assign w3015 = w2572 & w2881;
assign w3016 = w2842 | w2882;
assign w3017 = w2842 & w2882;
assign w3018 = w146 & w2883;
assign w3019 = w152 & w2884;
assign w3020 = w2567 & w2885;
assign w3021 = w2832 ~^ w2886;
assign w3022 = w2832 & w2887;
assign w3023 = w2851 ~^ w2889;
assign w3024 = w2851 | w2889;
assign w3025 = w2851 & w2889;
assign w3026 = w2835 ~^ w2891;
assign w3027 = w2835 & w2892;
assign w3028 = w152 & w2894;
assign w3029 = ~w2895;
assign w3030 = w145 & w2896;
assign w3031 = w149 & w2897;
assign w3032 = w2731 | w2898;
assign w3033 = ~w2899;
assign w3034 = w2790 ~^ w2900;
assign w3035 = w2790 ~| w2900;
assign w3036 = ~w2900;
assign w3037 = w2478 ~^ w2901;
assign w3038 = w2784 ~^ w2902;
assign w3039 = w2479 | w2903;
assign w3040 = w238 & w2904;
assign w3041 = w2608 & w2905;
assign w3042 = w2845 ~^ w2906;
assign w3043 = w231 & w2907;
assign w3044 = w2683 ~^ w2909;
assign w3045 = w237 & w2910;
assign w3046 = w2603 & w2911;
assign w3047 = ~w2915;
assign w3048 = w237 & w2916;
assign w3049 = w230 & w2918;
assign w3050 = w234 & w2919;
assign w3051 = w2760 | w2920;
assign w3052 = w2677 ~^ w2921;
assign w3053 = w2746 & w2923;
assign w3054 = w2899 ~^ w2924;
assign w3055 = ~w2924;
assign w3056 = w2751 & w2926;
assign w3057 = w2751 ~| w2926;
assign w3058 = w2504 ~^ w2927;
assign w3059 = w2504 & w2929;
assign w3060 = w2780 | w2930;
assign w3061 = w2438 ~| w2932;
assign w3062 = w2902 | w2934;
assign w3063 = w2925 | w2935;
assign w3064 = w347 & w2936;
assign w3065 = w2639 & w2937;
assign w3066 = w2845 | w2938;
assign w3067 = w2845 & w2938;
assign w3068 = w340 & w2939;
assign w3069 = w2826 ^ w2941;
assign w3070 = w346 & w2942;
assign w3071 = w2634 & w2943;
assign w3072 = w2912 | w2945;
assign w3073 = w346 & w2948;
assign w3074 = w339 & w2950;
assign w3075 = w343 & w2951;
assign w3076 = w2792 | w2952;
assign w3077 = w2806 | w2953;
assign w3078 = w2615 ~^ w2954;
assign w3079 = w2781 & w2954;
assign w3080 = ~w2956;
assign w3081 = w2956 ~^ w2957;
assign w3082 = w2697 ~^ w2959;
assign w3083 = w2858 & w2960;
assign w3084 = w2858 | w2960;
assign w3085 = w2818 | w2962;
assign w3086 = w2785 | w2963;
assign w3087 = w2859 ~^ w2964;
assign w3088 = w366 & w2965;
assign w3089 = w2675 & w2966;
assign w3090 = ~w2967;
assign w3091 = w359 & w2968;
assign w3092 = w2730 & w2970;
assign w3093 = w365 & w2971;
assign w3094 = w2670 & w2972;
assign w3095 = w2946 ~^ w2973;
assign w3096 = w2946 & w2973;
assign w3097 = w2946 ~| w2973;
assign w3098 = w2740 & w2974;
assign w3099 = w2914 ~^ w2975;
assign w3100 = w365 & w2977;
assign w3101 = ~w2978;
assign w3102 = w358 & w2979;
assign w3103 = w362 & w2980;
assign w3104 = w2827 | w2981;
assign w3105 = w2691 | w2983;
assign w3106 = w2949 & w2984;
assign w3107 = w2949 | w2984;
assign w3108 = w2848 | w2985;
assign w3109 = w2687 | w2987;
assign w3110 = ~w2989;
assign w3111 = ~w2990;
assign w3112 = w4 & w2991;
assign w3113 = w2816 | w2992;
assign w3114 = w2821 | w2993;
assign w3115 = w2712 | w2995;
assign w3116 = w2882 ~^ w2996;
assign w3117 = w2854 ~^ w2997;
assign w3118 = w2917 & w2997;
assign w3119 = w2917 | w2997;
assign w3120 = w2986 & w2998;
assign w3121 = w2986 | w2998;
assign w3122 = w2708 | w2999;
assign w3123 = w2453 ~| w3001;
assign w3124 = w1758 ~^ w3003;
assign w3125 = w2689 ~^ w3004;
assign w3126 = w2689 & w3004;
assign w3127 = w2689 | w3004;
assign w3128 = w2982 ~^ w3006;
assign w3129 = w2990 ~| w3007;
assign w3130 = ~w3007;
assign w3131 = w74 & w3008;
assign w3132 = w2874 | w3009;
assign w3133 = w2960 ~^ w3010;
assign w3134 = w2908 ~^ w3012;
assign w3135 = w2908 | w3012;
assign w3136 = w2908 & w3012;
assign w3137 = w2958 & w3013;
assign w3138 = ~w3014;
assign w3139 = w2738 | w3015;
assign w3140 = w2862 & w3016;
assign w3141 = w2870 ~^ w3018;
assign w3142 = ~w3018;
assign w3143 = w2998 ~^ w3019;
assign w3144 = w2734 | w3020;
assign w3145 = w2888 | w3022;
assign w3146 = w2913 ~^ w3023;
assign w3147 = w2913 & w3024;
assign w3148 = w2537 ~| w3027;
assign w3149 = w2994 ~^ w3030;
assign w3150 = w3007 ~^ w3031;
assign w3151 = ~w3031;
assign w3152 = w144 & w3032;
assign w3153 = w2877 ~^ w3034;
assign w3154 = w3011 | w3035;
assign w3155 = w2940 | w3036;
assign w3156 = w2820 | w3037;
assign w3157 = w2820 & w3037;
assign w3158 = w2776 ~^ w3038;
assign w3159 = w2961 & w3039;
assign w3160 = w3006 | w3040;
assign w3161 = w3006 & w3040;
assign w3162 = w2767 | w3041;
assign w3163 = w2938 ~^ w3042;
assign w3164 = w2978 ~^ w3043;
assign w3165 = ~w3043;
assign w3166 = ~w3045;
assign w3167 = w2763 | w3046;
assign w3168 = w2988 ~^ w3048;
assign w3169 = w2988 & w3048;
assign w3170 = w2988 | w3048;
assign w3171 = ~w3049;
assign w3172 = w229 & w3051;
assign w3173 = w2922 | w3053;
assign w3174 = w2967 ~^ w3054;
assign w3175 = ~w3054;
assign w3176 = w3033 | w3055;
assign w3177 = w2928 | w3059;
assign w3178 = w2704 ~^ w3060;
assign w3179 = ~w3060;
assign w3180 = w2933 | w3061;
assign w3181 = w3062 & w3063;
assign w3182 = w2989 ~| w3064;
assign w3183 = ~w3064;
assign w3184 = w2799 | w3065;
assign w3185 = w2906 & w3066;
assign w3186 = w2949 ~^ w3068;
assign w3187 = w3044 ^ w3069;
assign w3188 = ~w3070;
assign w3189 = w2795 | w3071;
assign w3190 = w3064 ~^ w3074;
assign w3191 = ~w3074;
assign w3192 = ~w3075;
assign w3193 = w338 & w3076;
assign w3194 = w2809 ~^ w3078;
assign w3195 = w2955 ~| w3078;
assign w3196 = ~w3078;
assign w3197 = w2749 | w3079;
assign w3198 = w2957 ~| w3080;
assign w3199 = w2957 & w3080;
assign w3200 = w2931 ~^ w3081;
assign w3201 = w3044 & w3082;
assign w3202 = w3044 ~| w3082;
assign w3203 = w2876 & w3084;
assign w3204 = w2704 ~| w3085;
assign w3205 = w2704 & w3085;
assign w3206 = w3058 ~^ w3087;
assign w3207 = w3058 & w3087;
assign w3208 = w3058 | w3087;
assign w3209 = w3049 ~^ w3088;
assign w3210 = ~w3088;
assign w3211 = w2834 | w3089;
assign w3212 = w3054 ~| w3090;
assign w3213 = w2870 ~| w3091;
assign w3214 = ~w3091;
assign w3215 = w2969 | w3092;
assign w3216 = w3070 ~^ w3093;
assign w3217 = ~w3093;
assign w3218 = w2830 | w3094;
assign w3219 = w3072 ~^ w3095;
assign w3220 = w3072 ~| w3097;
assign w3221 = ~w3099;
assign w3222 = w2944 ~^ w3100;
assign w3223 = ~w3100;
assign w3224 = w2994 | w3102;
assign w3225 = w2994 & w3102;
assign w3226 = w3075 ~^ w3103;
assign w3227 = ~w3103;
assign w3228 = w357 & w3104;
assign w3229 = w1 & w3105;
assign w3230 = w3068 & w3107;
assign w3231 = w8 & w3109;
assign w3232 = w3113 & w3114;
assign w3233 = w71 & w3115;
assign w3234 = ~w3116;
assign w3235 = w2917 ^ w3117;
assign w3236 = w2854 & w3119;
assign w3237 = w3019 & w3121;
assign w3238 = w78 & w3122;
assign w3239 = w3002 | w3123;
assign w3240 = w3028 ~^ w3125;
assign w3241 = w3028 & w3127;
assign w3242 = w3040 ~^ w3128;
assign w3243 = w3111 | w3130;
assign w3244 = w3112 & w3131;
assign w3245 = w3112 | w3131;
assign w3246 = ~w3133;
assign w3247 = w3052 ~^ w3134;
assign w3248 = w3052 & w3135;
assign w3249 = w2820 ~^ w3137;
assign w3250 = w141 & w3139;
assign w3251 = w3017 | w3140;
assign w3252 = w3091 ~^ w3141;
assign w3253 = w2986 ~^ w3143;
assign w3254 = w148 & w3144;
assign w3255 = w2564 ~^ w3145;
assign w3256 = w2564 & w3145;
assign w3257 = w2564 | w3145;
assign w3258 = ~w3146;
assign w3259 = w3025 | w3147;
assign w3260 = w3098 ~| w3148;
assign w3261 = w3102 ~^ w3149;
assign w3262 = w2990 ~^ w3150;
assign w3263 = w3129 | w3151;
assign w3264 = ~w3152;
assign w3265 = ~w3153;
assign w3266 = w3154 & w3155;
assign w3267 = w3137 | w3157;
assign w3268 = w2751 ~^ w3159;
assign w3269 = w3057 ~| w3159;
assign w3270 = w2982 & w3160;
assign w3271 = w226 & w3162;
assign w3272 = w3133 ~^ w3163;
assign w3273 = w3133 ~| w3163;
assign w3274 = ~w3163;
assign w3275 = w3101 | w3165;
assign w3276 = w233 & w3167;
assign w3277 = w3073 ~^ w3168;
assign w3278 = w3073 & w3170;
assign w3279 = w3045 ~^ w3172;
assign w3280 = ~w3172;
assign w3281 = w3108 ~^ w3174;
assign w3282 = w2967 | w3175;
assign w3283 = w2895 ~^ w3176;
assign w3284 = w3029 | w3176;
assign w3285 = ~w3176;
assign w3286 = w3085 ~^ w3178;
assign w3287 = w3158 ~^ w3180;
assign w3288 = ~w3180;
assign w3289 = w3110 | w3183;
assign w3290 = w335 & w3184;
assign w3291 = w3067 | w3185;
assign w3292 = w2984 ~^ w3186;
assign w3293 = w3082 ~^ w3187;
assign w3294 = w342 & w3189;
assign w3295 = w2989 ^ w3190;
assign w3296 = w3182 | w3191;
assign w3297 = w3045 ~| w3193;
assign w3298 = ~w3193;
assign out1[2] = w3077 ^ w3194;
assign w3299 = w2809 | w3196;
assign w3300 = w2931 ~| w3199;
assign w3301 = w3197 ~^ w3200;
assign w3302 = w3197 & w3200;
assign w3303 = w3197 | w3200;
assign w3304 = w3069 ~| w3202;
assign w3305 = w3083 | w3203;
assign w3306 = w3179 ~| w3204;
assign w3307 = w3086 ~^ w3206;
assign w3308 = w3086 & w3208;
assign w3309 = w3014 ~^ w3209;
assign w3310 = w3138 | w3209;
assign w3311 = ~w3209;
assign w3312 = w3171 | w3210;
assign w3313 = w354 & w3211;
assign w3314 = w3142 | w3213;
assign w3315 = w3005 | w3214;
assign w3316 = w3132 ~^ w3215;
assign w3317 = w3132 & w3215;
assign w3318 = w3132 | w3215;
assign w3319 = w3152 ~^ w3216;
assign w3320 = w3188 | w3217;
assign w3321 = w361 & w3218;
assign w3322 = ~w3219;
assign w3323 = w3096 | w3220;
assign w3324 = w3030 & w3224;
assign w3325 = w3192 | w3227;
assign w3326 = w3131 ~^ w3228;
assign w3327 = w3106 | w3230;
assign w3328 = w2868 ~^ w3231;
assign w3329 = w2868 | w3231;
assign w3330 = w2868 & w3231;
assign w3331 = w3177 ^ w3232;
assign w3332 = w3229 & w3233;
assign w3333 = w3229 | w3233;
assign w3334 = w3118 | w3236;
assign w3335 = w3120 | w3237;
assign w3336 = w2893 ~^ w3238;
assign w3337 = w2893 | w3238;
assign w3338 = w2893 & w3238;
assign w3339 = w3126 | w3241;
assign w3340 = w3228 & w3245;
assign w3341 = w3136 | w3248;
assign w3342 = w3037 ~^ w3249;
assign w3343 = w3226 ~^ w3250;
assign w3344 = ~w3250;
assign w3345 = ~w3251;
assign w3346 = ~w3254;
assign w3347 = w2890 ~^ w3259;
assign w3348 = w2739 | w3259;
assign w3349 = w2739 & w3259;
assign w3350 = w3124 ~^ w3260;
assign w3351 = w3242 & w3261;
assign w3352 = w3242 ~| w3261;
assign w3353 = ~w3262;
assign w3354 = w3243 & w3263;
assign w3355 = w3181 ~^ w3265;
assign w3356 = w3247 ^ w3266;
assign w3357 = w3156 & w3267;
assign w3358 = w2926 ~^ w3268;
assign w3359 = w3056 | w3269;
assign w3360 = w3161 | w3270;
assign w3361 = w3050 ~^ w3271;
assign w3362 = w3246 | w3274;
assign w3363 = ~w3277;
assign w3364 = w3169 | w3278;
assign w3365 = w3193 ~^ w3279;
assign w3366 = w3116 ~^ w3281;
assign w3367 = w3234 ~| w3281;
assign w3368 = ~w3281;
assign w3369 = w3108 & w3282;
assign w3370 = w3164 ~^ w3283;
assign w3371 = w2895 ~| w3285;
assign w3372 = w3177 & w3286;
assign w3373 = w3177 ~| w3286;
assign w3374 = w3158 ~| w3288;
assign w3375 = w3158 & w3288;
assign w3376 = w3050 | w3290;
assign w3377 = w3050 & w3290;
assign w3378 = ~w3291;
assign w3379 = w3235 ^ w3292;
assign w3380 = w3252 ~| w3292;
assign w3381 = w3252 & w3292;
assign w3382 = w3247 & w3293;
assign w3383 = w3247 ~| w3293;
assign w3384 = w2947 ~^ w3294;
assign w3385 = w2852 | w3294;
assign w3386 = w2852 & w3294;
assign w3387 = w3242 ^ w3295;
assign w3388 = w3289 & w3296;
assign w3389 = w3280 | w3297;
assign w3390 = w3166 | w3298;
assign w3391 = w3077 & w3299;
assign w3392 = w3198 | w3300;
assign w3393 = w3201 | w3304;
assign w3394 = w3251 ~^ w3305;
assign w3395 = w3251 ~| w3305;
assign w3396 = ~w3305;
assign w3397 = w3205 | w3306;
assign w3398 = w3153 ~| w3307;
assign w3399 = ~w3307;
assign w3400 = w3207 | w3308;
assign w3401 = w3275 ~^ w3309;
assign w3402 = w3014 ~| w3311;
assign w3403 = ~w3312;
assign w3404 = w3233 ~^ w3313;
assign w3405 = w3314 & w3315;
assign w3406 = w3173 ~^ w3316;
assign w3407 = w3173 & w3318;
assign w3408 = w2915 ~^ w3321;
assign w3409 = ~w3321;
assign w3410 = w3239 ~^ w3323;
assign w3411 = w3239 | w3323;
assign w3412 = w3239 & w3323;
assign w3413 = w3225 | w3324;
assign w3414 = w3319 ~^ w3325;
assign w3415 = w3264 ~| w3325;
assign w3416 = w3264 & w3325;
assign w3417 = w3112 ~^ w3326;
assign w3418 = ~w3327;
assign w3419 = w3276 ~^ w3328;
assign w3420 = w3276 & w3329;
assign w3421 = w3286 ~^ w3331;
assign w3422 = w3313 & w3333;
assign w3423 = w3327 ~| w3334;
assign w3424 = ~w3334;
assign w3425 = ~w3335;
assign w3426 = w2976 ~^ w3336;
assign w3427 = w2976 & w3337;
assign w3428 = w3146 ~^ w3339;
assign w3429 = w3146 ~| w3339;
assign w3430 = ~w3339;
assign w3431 = w3244 | w3340;
assign w3432 = w3287 ~^ w3342;
assign w3433 = w3312 ~^ w3343;
assign w3434 = w3312 | w3344;
assign w3435 = w3320 ~| w3346;
assign w3436 = w3320 & w3346;
assign w3437 = w1411 & w3348;
assign w3438 = w3295 ~| w3352;
assign w3439 = w3307 ~^ w3355;
assign w3440 = w3293 ^ w3356;
assign w3441 = w3357 ~^ w3358;
assign w3442 = ~w3358;
assign w3443 = ~w3359;
assign w3444 = w3290 ~^ w3361;
assign w3445 = w3255 ~^ w3364;
assign w3446 = w3257 & w3364;
assign w3447 = w3116 | w3368;
assign w3448 = w3212 | w3369;
assign w3449 = w3164 | w3371;
assign w3450 = w3232 ~| w3373;
assign w3451 = w3342 ~| w3375;
assign w3452 = w3271 & w3376;
assign w3453 = w3252 ~^ w3379;
assign w3454 = w3235 ~| w3380;
assign w3455 = w3266 ~| w3383;
assign w3456 = w2852 ~^ w3384;
assign w3457 = w2947 & w3385;
assign w3458 = w3261 ~^ w3387;
assign w3459 = w3389 & w3390;
assign w3460 = w3195 | w3391;
assign w3461 = w3366 ~^ w3393;
assign w3462 = w3291 ~^ w3394;
assign w3463 = w3378 | w3395;
assign w3464 = w3345 | w3396;
assign w3465 = w3272 ~^ w3397;
assign w3466 = ~w3397;
assign w3467 = w3181 | w3398;
assign w3468 = w3265 | w3399;
assign w3469 = ~w3401;
assign w3470 = w3275 | w3402;
assign w3471 = w3250 ~| w3403;
assign w3472 = w3229 ~^ w3404;
assign w3473 = w3334 ^ w3405;
assign w3474 = w3341 ~^ w3406;
assign w3475 = w3341 | w3406;
assign w3476 = w3341 & w3406;
assign w3477 = w3317 | w3407;
assign w3478 = w3254 ~^ w3408;
assign w3479 = w3047 | w3409;
assign w3480 = w3347 ~^ w3410;
assign w3481 = w3347 & w3411;
assign w3482 = w3388 ^ w3413;
assign w3483 = w3360 ~| w3413;
assign w3484 = w3360 & w3413;
assign w3485 = w3365 ~^ w3414;
assign w3486 = w3365 | w3414;
assign w3487 = w3365 & w3414;
assign w3488 = w3216 ~| w3416;
assign w3489 = ~w3417;
assign w3490 = w3330 | w3420;
assign w3491 = w3359 | w3421;
assign w3492 = ~w3421;
assign w3493 = w3332 | w3422;
assign w3494 = w3405 | w3423;
assign w3495 = w3418 | w3424;
assign w3496 = w3419 ~^ w3426;
assign w3497 = w3419 & w3426;
assign w3498 = w3419 | w3426;
assign w3499 = w3338 | w3427;
assign w3500 = w3000 ~^ w3428;
assign w3501 = w3000 | w3429;
assign w3502 = w3258 | w3430;
assign w3503 = w3392 ~^ w3432;
assign w3504 = w3392 & w3432;
assign w3505 = w3392 | w3432;
assign w3506 = w3408 ~| w3436;
assign w3507 = w3349 | w3437;
assign w3508 = w3351 | w3438;
assign w3509 = w3439 ~^ w3441;
assign w3510 = w3439 & w3442;
assign w3511 = w3439 ~| w3442;
assign w3512 = w3421 ~^ w3443;
assign w3513 = w3433 & w3444;
assign w3514 = w3433 ~| w3444;
assign w3515 = ~w3445;
assign w3516 = w3256 | w3446;
assign w3517 = w3393 & w3447;
assign w3518 = w3370 | w3448;
assign w3519 = w3370 & w3448;
assign w3520 = w3284 & w3449;
assign w3521 = w3372 | w3450;
assign w3522 = w3374 | w3451;
assign w3523 = w3377 | w3452;
assign w3524 = w3381 | w3454;
assign w3525 = w3382 | w3455;
assign w3526 = w3335 ~| w3456;
assign w3527 = ~w3456;
assign w3528 = w3386 | w3457;
assign w3529 = w3425 ~^ w3459;
assign out1[3] = w3301 ~^ w3460;
assign w3530 = w3303 & w3460;
assign w3531 = ~w3461;
assign w3532 = w3453 & w3462;
assign w3533 = w3453 ~| w3462;
assign w3534 = w3463 & w3464;
assign w3535 = w3461 ~^ w3465;
assign w3536 = ~w3465;
assign w3537 = w3273 | w3466;
assign w3538 = w3467 & w3468;
assign w3539 = w3310 & w3470;
assign w3540 = w3226 | w3471;
assign w3541 = w3262 ~^ w3472;
assign w3542 = w3262 ~| w3472;
assign w3543 = ~w3472;
assign w3544 = w3327 ~^ w3473;
assign w3545 = w3448 ~^ w3477;
assign w3546 = w3320 ~^ w3478;
assign w3547 = w3222 ~^ w3479;
assign w3548 = w3223 ~| w3479;
assign w3549 = w3223 & w3479;
assign w3550 = w3412 | w3481;
assign w3551 = w3360 ~^ w3482;
assign w3552 = w3388 ~| w3483;
assign w3553 = w3415 | w3488;
assign w3554 = w3277 ~^ w3490;
assign w3555 = w3240 & w3490;
assign w3556 = w3240 ~| w3490;
assign w3557 = w3400 & w3491;
assign w3558 = w3443 ~| w3492;
assign w3559 = w3253 ~| w3493;
assign w3560 = w3253 & w3493;
assign w3561 = w3354 ^ w3493;
assign w3562 = w3494 & w3495;
assign w3563 = w3431 ~^ w3496;
assign w3564 = w3431 & w3498;
assign w3565 = w3021 ~^ w3499;
assign w3566 = ~w3500;
assign w3567 = w3501 & w3502;
assign w3568 = w3435 | w3506;
assign w3569 = w3350 ~^ w3507;
assign w3570 = ~w3508;
assign w3571 = w3357 ~| w3511;
assign w3572 = w3400 ~^ w3512;
assign w3573 = w3026 ~^ w3516;
assign w3574 = w3367 | w3517;
assign w3575 = w3477 & w3518;
assign w3576 = w3469 & w3520;
assign w3577 = w3469 ~| w3520;
assign w3578 = w3474 ~^ w3521;
assign w3579 = w3475 & w3521;
assign w3580 = w3509 ~^ w3522;
assign w3581 = w3509 & w3522;
assign w3582 = w3509 | w3522;
assign w3583 = w3417 ~^ w3523;
assign w3584 = w3417 ~| w3523;
assign w3585 = ~w3523;
assign w3586 = ~w3525;
assign w3587 = w3459 | w3526;
assign w3588 = w3425 | w3527;
assign w3589 = w3499 | w3528;
assign w3590 = w3499 & w3528;
assign w3591 = w3456 ~^ w3529;
assign w3592 = w3302 | w3530;
assign w3593 = w3465 ~| w3531;
assign w3594 = w3520 ~^ w3534;
assign w3595 = w3525 ~^ w3535;
assign w3596 = w3461 | w3536;
assign w3597 = w3362 & w3537;
assign w3598 = w3440 ^ w3538;
assign w3599 = w3434 & w3540;
assign w3600 = w3539 ^ w3541;
assign w3601 = w3539 | w3542;
assign w3602 = w3353 | w3543;
assign w3603 = w3524 ~^ w3544;
assign w3604 = w3524 | w3544;
assign w3605 = w3524 & w3544;
assign w3606 = w3370 ~^ w3545;
assign w3607 = ~w3546;
assign w3608 = ~w3547;
assign w3609 = w2944 ~| w3549;
assign w3610 = w3221 ~^ w3550;
assign w3611 = w3508 ~^ w3551;
assign w3612 = w3508 ~| w3551;
assign w3613 = ~w3551;
assign w3614 = w3484 | w3552;
assign w3615 = w3546 | w3553;
assign w3616 = ~w3553;
assign w3617 = w3240 ~^ w3554;
assign w3618 = w3363 ~| w3556;
assign w3619 = w3557 | w3558;
assign w3620 = w3354 ~| w3559;
assign w3621 = w3253 ^ w3561;
assign w3622 = w3514 ~| w3562;
assign w3623 = w3444 ^ w3562;
assign w3624 = w3497 | w3564;
assign w3625 = w3528 ~^ w3565;
assign w3626 = ~w3567;
assign w3627 = w3547 ~^ w3568;
assign w3628 = w3547 ~| w3568;
assign w3629 = ~w3568;
assign w3630 = w3510 | w3571;
assign w3631 = w3440 | w3572;
assign w3632 = w3440 & w3572;
assign w3633 = w3567 ~^ w3573;
assign w3634 = w3519 | w3575;
assign w3635 = w3534 ~| w3576;
assign w3636 = ~w3578;
assign w3637 = w3476 | w3579;
assign w3638 = w3489 | w3585;
assign w3639 = w3587 & w3588;
assign w3640 = w3021 & w3589;
assign w3641 = w3563 & w3591;
assign w3642 = w3563 ~| w3591;
assign out1[4] = w3503 ~^ w3592;
assign w3643 = w3505 & w3592;
assign w3644 = w3586 | w3593;
assign w3645 = w3401 ~^ w3594;
assign w3646 = ~w3595;
assign w3647 = w3533 ~| w3597;
assign w3648 = w3462 ^ w3597;
assign w3649 = w3572 ~^ w3598;
assign w3650 = w3583 ~^ w3599;
assign w3651 = w3584 | w3599;
assign w3652 = ~w3600;
assign w3653 = w3601 & w3602;
assign w3654 = w3574 ~^ w3606;
assign w3655 = w3574 | w3606;
assign w3656 = w3574 & w3606;
assign w3657 = w3548 | w3609;
assign w3658 = w3600 ~^ w3611;
assign w3659 = w3570 | w3613;
assign w3660 = w3485 ~^ w3614;
assign w3661 = w3486 & w3614;
assign w3662 = w3546 ~^ w3616;
assign w3663 = w3607 ~| w3616;
assign w3664 = w3555 | w3618;
assign w3665 = w3578 ~^ w3619;
assign w3666 = w3560 | w3620;
assign w3667 = w3513 | w3622;
assign w3668 = w3433 ~^ w3623;
assign w3669 = ~w3624;
assign w3670 = w3617 & w3625;
assign w3671 = w3617 ~| w3625;
assign w3672 = w3516 | w3626;
assign w3673 = w3516 & w3626;
assign w3674 = w3624 ~^ w3627;
assign w3675 = w3608 | w3629;
assign w3676 = w3538 | w3632;
assign w3677 = w3603 ~^ w3634;
assign w3678 = w3604 & w3634;
assign w3679 = w3577 | w3635;
assign w3680 = w3595 ~| w3636;
assign w3681 = w3625 ^ w3639;
assign w3682 = w3590 | w3640;
assign w3683 = w3504 | w3643;
assign w3684 = w3596 & w3644;
assign w3685 = w3458 ~^ w3645;
assign w3686 = w3458 | w3645;
assign w3687 = w3458 & w3645;
assign w3688 = w3578 | w3646;
assign w3689 = w3532 | w3647;
assign w3690 = w3453 ~^ w3648;
assign w3691 = w3630 ~^ w3649;
assign w3692 = w3630 | w3649;
assign w3693 = w3630 & w3649;
assign w3694 = w3621 ~| w3650;
assign w3695 = w3621 & w3650;
assign w3696 = w3638 & w3651;
assign w3697 = w3612 | w3652;
assign w3698 = w3621 ^ w3653;
assign w3699 = w3637 ~^ w3654;
assign w3700 = w3637 & w3655;
assign w3701 = w3219 ~^ w3657;
assign w3702 = w3322 ~| w3657;
assign w3703 = ~w3657;
assign w3704 = ~w3658;
assign w3705 = w3487 | w3661;
assign w3706 = w3566 | w3664;
assign w3707 = ~w3664;
assign w3708 = w3595 ~^ w3665;
assign w3709 = w3662 ~^ w3666;
assign w3710 = w3615 & w3666;
assign w3711 = w3660 ~^ w3667;
assign w3712 = w3660 | w3667;
assign w3713 = w3660 & w3667;
assign w3714 = w3628 | w3669;
assign w3715 = w3639 ~| w3671;
assign w3716 = w3026 & w3672;
assign w3717 = ~w3674;
assign w3718 = w3631 & w3676;
assign w3719 = w3605 | w3678;
assign w3720 = w3668 ~^ w3679;
assign w3721 = w3668 & w3679;
assign w3722 = w3668 | w3679;
assign w3723 = w3617 ~^ w3681;
assign w3724 = w3664 ~^ w3682;
assign out1[5] = w3580 ~^ w3683;
assign w3725 = w3582 & w3683;
assign w3726 = w3619 & w3688;
assign w3727 = w3685 ~^ w3689;
assign w3728 = w3686 & w3689;
assign w3729 = w3684 ^ w3690;
assign w3730 = w3653 ~| w3695;
assign w3731 = w3642 ~| w3696;
assign w3732 = w3591 ^ w3696;
assign w3733 = w3659 & w3697;
assign w3734 = w3650 ~^ w3698;
assign w3735 = w3690 & w3699;
assign w3736 = w3690 ~| w3699;
assign w3737 = w3656 | w3700;
assign w3738 = w3445 ~^ w3701;
assign w3739 = w3515 | w3702;
assign w3740 = w3219 | w3703;
assign w3741 = w3682 & w3706;
assign w3742 = w3500 ~| w3707;
assign w3743 = w3705 ~^ w3709;
assign w3744 = ~w3709;
assign w3745 = w3663 | w3710;
assign w3746 = w3675 & w3714;
assign w3747 = w3670 | w3715;
assign w3748 = w3673 | w3716;
assign w3749 = w3708 ~^ w3718;
assign w3750 = w3708 | w3718;
assign w3751 = w3708 & w3718;
assign w3752 = w3719 ~^ w3720;
assign w3753 = w3719 & w3722;
assign w3754 = w3500 ~^ w3724;
assign w3755 = w3581 | w3725;
assign w3756 = w3680 | w3726;
assign w3757 = w3677 ~^ w3727;
assign w3758 = w3677 & w3727;
assign w3759 = w3677 | w3727;
assign w3760 = w3687 | w3728;
assign w3761 = w3699 ~^ w3729;
assign w3762 = w3694 | w3730;
assign w3763 = w3641 | w3731;
assign w3764 = w3563 ~^ w3732;
assign w3765 = ~w3733;
assign w3766 = w3711 ~^ w3734;
assign w3767 = w3712 & w3734;
assign w3768 = w3684 ~| w3736;
assign w3769 = w3739 & w3740;
assign w3770 = w3741 | w3742;
assign w3771 = w3705 | w3744;
assign w3772 = w3705 & w3744;
assign w3773 = w3717 ~^ w3745;
assign w3774 = w3674 | w3745;
assign w3775 = ~w3745;
assign w3776 = w3738 ~^ w3746;
assign w3777 = w3610 ~^ w3748;
assign w3778 = w3704 ~^ w3752;
assign w3779 = w3658 | w3752;
assign w3780 = ~w3752;
assign w3781 = w3721 | w3753;
assign w3782 = w3746 | w3754;
assign w3783 = w3746 & w3754;
assign out1[6] = w3691 ~^ w3755;
assign w3784 = w3692 & w3755;
assign w3785 = ~w3756;
assign w3786 = w3737 ~^ w3757;
assign w3787 = w3737 & w3759;
assign w3788 = w3756 ~^ w3761;
assign w3789 = w3756 ~| w3761;
assign w3790 = ~w3761;
assign w3791 = w3743 ~^ w3762;
assign w3792 = ~w3763;
assign w3793 = ~w3764;
assign w3794 = w3765 | w3766;
assign w3795 = ~w3766;
assign w3796 = w3713 | w3767;
assign w3797 = w3735 | w3768;
assign w3798 = w3480 ^ w3769;
assign w3799 = w3480 ~| w3770;
assign w3800 = w3480 & w3770;
assign w3801 = w3762 & w3771;
assign w3802 = w3723 ~^ w3773;
assign w3803 = w3723 & w3774;
assign w3804 = w3717 ~| w3775;
assign w3805 = w3754 ~^ w3776;
assign w3806 = w3569 ~^ w3777;
assign w3807 = w3760 ~^ w3778;
assign w3808 = w3760 & w3779;
assign w3809 = w3704 ~| w3780;
assign w3810 = w3765 ~^ w3781;
assign w3811 = w3738 | w3783;
assign w3812 = w3693 | w3784;
assign w3813 = ~w3786;
assign w3814 = w3758 | w3787;
assign w3815 = w3785 | w3790;
assign w3816 = ~w3791;
assign w3817 = w3791 ~| w3793;
assign w3818 = w3781 & w3794;
assign w3819 = w3733 ~| w3795;
assign w3820 = w3786 ~| w3797;
assign w3821 = ~w3797;
assign w3822 = w3770 ~^ w3798;
assign w3823 = w3769 ~| w3799;
assign w3824 = w3772 | w3801;
assign w3825 = w3792 | w3802;
assign w3826 = ~w3802;
assign w3827 = w3803 | w3804;
assign w3828 = w3747 ^ w3805;
assign w3829 = w3808 | w3809;
assign w3830 = w3795 ~^ w3810;
assign w3831 = w3782 & w3811;
assign out1[7] = w3749 ~^ w3812;
assign w3832 = ~w3812;
assign w3833 = w3797 ~^ w3813;
assign w3834 = w3807 ~^ w3814;
assign w3835 = ~w3814;
assign w3836 = w3793 ~^ w3816;
assign w3837 = w3764 | w3816;
assign w3838 = w3818 | w3819;
assign w3839 = w3813 | w3821;
assign w3840 = w3633 ~^ w3822;
assign w3841 = ~w3822;
assign w3842 = w3800 ~| w3823;
assign w3843 = ~w3824;
assign w3844 = w3792 ~^ w3826;
assign w3845 = w3763 ~| w3826;
assign w3846 = w3747 ~| w3827;
assign w3847 = w3747 & w3827;
assign w3848 = w3827 ~^ w3828;
assign w3849 = ~w3829;
assign w3850 = ~w3830;
assign w3851 = w3633 ~| w3831;
assign w3852 = w3633 & w3831;
assign w3853 = w3751 | w3832;
assign w3854 = w3807 & w3835;
assign w3855 = w3807 ~| w3835;
assign w3856 = w3796 ~^ w3836;
assign w3857 = w3796 & w3837;
assign w3858 = ~w3838;
assign w3859 = w3831 ~^ w3840;
assign w3860 = w3806 ~^ w3842;
assign w3861 = w3824 ~^ w3844;
assign w3862 = w3843 | w3845;
assign w3863 = w3805 ~| w3846;
assign w3864 = ~w3848;
assign w3865 = w3830 | w3849;
assign w3866 = w3829 ~^ w3850;
assign w3867 = w3829 ~| w3850;
assign w3868 = w3841 ~| w3852;
assign w3869 = w3750 & w3853;
assign w3870 = w3838 ~^ w3856;
assign w3871 = w3817 | w3857;
assign w3872 = w3856 ~| w3858;
assign w3873 = w3856 & w3858;
assign w3874 = ~w3861;
assign w3875 = w3825 & w3862;
assign w3876 = w3847 | w3863;
assign w3877 = w3851 ~| w3868;
assign w3878 = w3789 | w3869;
assign out1[8] = w3788 ^ w3869;
assign w3879 = ~w3871;
assign w3880 = w3871 ~^ w3874;
assign w3881 = w3871 ~| w3874;
assign w3882 = w3848 ~^ w3875;
assign w3883 = w3864 & w3875;
assign w3884 = w3864 ~| w3875;
assign w3885 = w3859 ~^ w3876;
assign w3886 = w3859 | w3876;
assign w3887 = w3859 & w3876;
assign w3888 = w3860 ~^ w3877;
assign w3889 = w3815 & w3878;
assign w3890 = w3861 | w3879;
assign out1[9] = w3833 ~^ w3889;
assign w3891 = w3820 | w3889;
assign w3892 = w3839 & w3891;
assign out1[10] = w3834 ~^ w3892;
assign w3893 = w3854 ~| w3892;
assign w3894 = w3855 | w3893;
assign out1[11] = w3866 ~^ w3894;
assign w3895 = ~w3894;
assign w3896 = w3867 | w3895;
assign w3897 = w3865 & w3896;
assign out1[12] = w3870 ~^ w3897;
assign w3898 = w3873 ~| w3897;
assign w3899 = w3872 | w3898;
assign out1[13] = w3880 ~^ w3899;
assign w3900 = ~w3899;
assign w3901 = w3881 | w3900;
assign w3902 = w3890 & w3901;
assign out1[14] = w3882 ~^ w3902;
assign w3903 = w3883 ~| w3902;
assign w3904 = w3884 | w3903;
assign out1[15] = w3885 ~^ w3904;
assign w3905 = w3886 & w3904;
assign w3906 = w3887 ~| w3905;
assign out1[16] = w3888 ~^ w3906;
wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906;
endmodule
module top(in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, out1, out2, out3);
input wire [12:0] in1;
input wire [17:0] in2;
input wire [31:0] in3;
input wire [31:0] in7;
input wire [31:0] in9;
input wire in4;
input wire in5;
input wire in6;
input wire in8;
input wire [4:0] in10;
input wire [15:0] in11;
output wire [32:0] out1;
output wire [31:0] out2;
output wire [31:0] out3;
assign w0 = ~in1[0];
assign w1 = ~in1[0];
assign w2 = ~in1[0];
assign w3 = ~in1[0];
assign w4 = ~in1[0];
assign w5 = ~in1[0];
assign w6 = ~in1[0];
assign w7 = ~in1[0];
assign w8 = ~in1[0];
assign w9 = ~in1[1];
assign w10 = in1[1] & in1[0];
assign w11 = ~in1[1];
assign w12 = ~in1[1];
assign w13 = ~in1[2];
assign w14 = in1[2] ~| in1[1];
assign w15 = ~in1[2];
assign w16 = ~in1[3];
assign w17 = in1[3] ~^ in1[2];
assign w18 = ~in1[3];
assign w19 = ~in1[4];
assign w20 = in1[4] ~| in1[3];
assign w21 = ~in1[4];
assign w22 = ~in1[5];
assign w23 = in1[5] ~^ in1[4];
assign w24 = ~in1[5];
assign w25 = ~in1[6];
assign w26 = in1[6] ~| in1[5];
assign w27 = ~in1[6];
assign w28 = ~in1[7];
assign w29 = in1[7] ~^ in1[6];
assign w30 = ~in1[7];
assign w31 = ~in1[8];
assign w32 = in1[8] ~| in1[7];
assign w33 = ~in1[8];
assign w34 = ~in1[9];
assign w35 = in1[9] ~^ in1[8];
assign w36 = ~in1[9];
assign w37 = ~in1[10];
assign w38 = in1[10] ~| in1[9];
assign w39 = ~in1[10];
assign w40 = ~in1[11];
assign w41 = in1[11] ~^ in1[10];
assign w42 = ~in1[11];
assign w43 = ~in1[12];
assign w44 = in1[12] ~^ in1[11];
assign w45 = ~in1[12];
assign w46 = in1[7] ~^ in2[1];
assign w47 = in1[3] ~^ in2[1];
assign w48 = in1[9] ~^ in2[1];
assign w49 = in1[5] ~^ in2[1];
assign w50 = in1[1] ~^ in2[1];
assign w51 = in1[11] ~^ in2[1];
assign w52 = in1[5] ~^ in2[2];
assign w53 = in1[3] ~^ in2[2];
assign w54 = in1[9] ~^ in2[2];
assign w55 = in1[7] ~^ in2[2];
assign w56 = in1[1] ~^ in2[2];
assign w57 = in1[11] ~^ in2[2];
assign w58 = in1[9] ~^ in2[3];
assign w59 = in1[5] ~^ in2[3];
assign w60 = in1[3] ~^ in2[3];
assign w61 = in1[7] ~^ in2[3];
assign w62 = in1[1] ~^ in2[3];
assign w63 = in1[11] ~^ in2[3];
assign w64 = in1[5] ~^ in2[4];
assign w65 = in1[7] ~^ in2[4];
assign w66 = in1[3] ~^ in2[4];
assign w67 = in1[9] ~^ in2[4];
assign w68 = in1[1] ~^ in2[4];
assign w69 = in1[11] ~^ in2[4];
assign w70 = in1[5] ~^ in2[5];
assign w71 = in1[9] ~^ in2[5];
assign w72 = in1[7] ~^ in2[5];
assign w73 = in1[3] ~^ in2[5];
assign w74 = in1[1] ~^ in2[5];
assign w75 = in1[11] ~^ in2[5];
assign w76 = in1[9] ~^ in2[6];
assign w77 = in1[7] ~^ in2[6];
assign w78 = in1[5] ~^ in2[6];
assign w79 = in1[3] ~^ in2[6];
assign w80 = in1[1] ~^ in2[6];
assign w81 = in1[11] ~^ in2[6];
assign w82 = in1[9] ~^ in2[7];
assign w83 = in1[7] ~^ in2[7];
assign w84 = in1[5] ~^ in2[7];
assign w85 = in1[3] ~^ in2[7];
assign w86 = in1[1] ~^ in2[7];
assign w87 = in1[11] ~^ in2[7];
assign w88 = ~in2[7];
assign w89 = in1[9] ~^ in2[8];
assign w90 = in1[5] ~^ in2[8];
assign w91 = in1[3] ~^ in2[8];
assign w92 = in1[7] ~^ in2[8];
assign w93 = in1[1] ~^ in2[8];
assign w94 = in1[11] ~^ in2[8];
assign w95 = ~in2[8];
assign w96 = in1[7] ~^ in2[9];
assign w97 = in1[3] ~^ in2[9];
assign w98 = in1[9] ~^ in2[9];
assign w99 = in1[5] ~^ in2[9];
assign w100 = in1[1] ~^ in2[9];
assign w101 = in1[11] ~^ in2[9];
assign w102 = in1[5] ~^ in2[10];
assign w103 = in1[3] ~^ in2[10];
assign w104 = in1[9] ~^ in2[10];
assign w105 = in1[1] ~^ in2[10];
assign w106 = in1[7] ~^ in2[10];
assign w107 = in1[11] ~^ in2[10];
assign w108 = in1[3] ~^ in2[11];
assign w109 = in1[9] ~^ in2[11];
assign w110 = in1[7] ~^ in2[11];
assign w111 = in1[5] ~^ in2[11];
assign w112 = in1[1] ~^ in2[11];
assign w113 = in1[11] ~^ in2[11];
assign w114 = in1[5] ~^ in2[12];
assign w115 = in1[9] ~^ in2[12];
assign w116 = in1[7] ~^ in2[12];
assign w117 = in1[3] ~^ in2[12];
assign w118 = in1[1] ~^ in2[12];
assign w119 = in1[11] ~^ in2[12];
assign w120 = in1[7] ~^ in2[13];
assign w121 = in1[9] ~^ in2[13];
assign w122 = in1[3] ~^ in2[13];
assign w123 = in1[1] ~^ in2[13];
assign w124 = in1[5] ~^ in2[13];
assign w125 = in1[11] ~^ in2[13];
assign w126 = in1[9] ~^ in2[14];
assign w127 = in1[5] ~^ in2[14];
assign w128 = in1[3] ~^ in2[14];
assign w129 = in1[7] ~^ in2[14];
assign w130 = in1[1] ~^ in2[14];
assign w131 = in1[11] ~^ in2[14];
assign w132 = in1[9] ~^ in2[15];
assign w133 = in1[5] ~^ in2[15];
assign w134 = in1[7] ~^ in2[15];
assign w135 = in1[3] ~^ in2[15];
assign w136 = in1[1] ~^ in2[15];
assign w137 = in1[11] ~^ in2[15];
assign w138 = in1[5] ~^ in2[16];
assign w139 = in1[7] ~^ in2[16];
assign w140 = in1[3] ~^ in2[16];
assign w141 = in1[9] ~^ in2[16];
assign w142 = in1[1] ~^ in2[16];
assign w143 = in1[11] ~^ in2[16];
assign w144 = in1[9] ~^ in2[17];
assign w145 = in1[5] ~^ in2[17];
assign w146 = in1[3] ~^ in2[17];
assign w147 = in1[7] ~^ in2[17];
assign w148 = in1[1] ~^ in2[17];
assign w149 = in1[11] ~^ in2[17];
assign w150 = ~in2[17];
assign w151 = ~in3[0];
assign w152 = ~in3[1];
assign w153 = ~in3[2];
assign w154 = ~in3[3];
assign w155 = ~in3[4];
assign w156 = ~in3[5];
assign w157 = ~in3[6];
assign w158 = ~in3[7];
assign w159 = ~in3[8];
assign w160 = ~in3[9];
assign w161 = ~in3[10];
assign w162 = ~in3[11];
assign w163 = ~in3[12];
assign w164 = ~in3[17];
assign w165 = ~in3[18];
assign w166 = ~in3[19];
assign w167 = ~in3[20];
assign w168 = in3[21] ~^ in3[20];
assign w169 = in3[21] ~| in3[20];
assign w170 = ~in3[21];
assign w171 = ~in3[22];
assign w172 = in3[23] ~^ in3[22];
assign w173 = in3[23] ~| in3[22];
assign w174 = ~in3[23];
assign w175 = ~in3[24];
assign w176 = in3[25] ~^ in3[24];
assign w177 = in3[25] ~| in3[24];
assign w178 = ~in3[25];
assign w179 = ~in3[26];
assign w180 = in3[27] ~^ in3[26];
assign w181 = in3[27] & in3[26];
assign w182 = in3[27] | in3[26];
assign w183 = ~in3[28];
assign w184 = in3[29] ~^ in3[28];
assign w185 = in3[29] ~| in3[28];
assign w186 = ~in3[29];
assign w187 = in3[31] ~^ in3[30];
assign w188 = in3[31] ~| in3[30];
assign w189 = ~in9[2];
assign w190 = ~in9[4];
assign w191 = ~in9[5];
assign w192 = ~in9[6];
assign w193 = ~in9[7];
assign w194 = ~in9[8];
assign w195 = ~in9[9];
assign w196 = ~in9[10];
assign w197 = ~in9[11];
assign w198 = ~in9[12];
assign w199 = ~in9[13];
assign w200 = ~in9[14];
assign w201 = ~in9[15];
assign w202 = ~in9[16];
assign w203 = ~in4;
assign w204 = ~in4;
assign w205 = ~in5;
assign w206 = ~in5;
assign w207 = ~in6;
assign w208 = ~in6;
assign w209 = ~in6;
assign w210 = ~in6;
assign w211 = ~in6;
assign w212 = ~in6;
assign w213 = ~in6;
assign w214 = ~in6;
assign w215 = ~in6;
assign w216 = ~in6;
assign w217 = ~in6;
assign w218 = ~in6;
assign w219 = ~in6;
assign w220 = ~in6;
assign w221 = ~in6;
assign w222 = in6 ~| in7[5];
assign w223 = in6 ~| in7[13];
assign w224 = in6 ~| in7[4];
assign w225 = in6 ~| in7[25];
assign w226 = in6 ~| in7[3];
assign w227 = in6 ~| in7[15];
assign w228 = in6 ~| in7[18];
assign w229 = in6 ~| in7[2];
assign w230 = in6 ~| in7[1];
assign w231 = in6 ~| in7[24];
assign w232 = in6 ~| in7[21];
assign w233 = in6 ~| in7[29];
assign w234 = in6 ~| in7[9];
assign w235 = in6 ~| in7[0];
assign w236 = in6 ~| in7[7];
assign w237 = in6 ~| in7[28];
assign w238 = ~in6;
assign w239 = ~in6;
assign w240 = ~in6;
assign w241 = ~in6;
assign w242 = ~in6;
assign w243 = ~in6;
assign w244 = ~in6;
assign w245 = ~in6;
assign w246 = in6 ~| in7[26];
assign w247 = in6 ~| in7[23];
assign w248 = in6 ~| in7[6];
assign w249 = in6 ~| in7[16];
assign w250 = in6 ~| in7[30];
assign w251 = in6 ~| in7[12];
assign w252 = in6 ~| in7[19];
assign w253 = in6 ~| in7[31];
assign w254 = in6 ~| in7[10];
assign w255 = in6 ~| in7[14];
assign w256 = in6 ~| in7[11];
assign w257 = in6 ~| in7[20];
assign w258 = in6 ~| in7[27];
assign w259 = in6 ~| in7[8];
assign w260 = in6 ~| in7[17];
assign w261 = in6 ~| in7[22];
assign w262 = in1[0] & in10[0];
assign w263 = in1[1] & in10[0];
assign w264 = ~in10[0];
assign w265 = ~in10[0];
assign w266 = ~in10[0];
assign w267 = ~in10[0];
assign w268 = ~in10[0];
assign w269 = ~in10[0];
assign w270 = ~in10[1];
assign w271 = ~in10[1];
assign w272 = ~in10[1];
assign w273 = ~in10[1];
assign w274 = ~in10[1];
assign w275 = ~in10[1];
assign w276 = in1[6] & in10[2];
assign w277 = in1[7] & in10[2];
assign w278 = in1[5] & in10[2];
assign w279 = ~in10[2];
assign w280 = ~in10[2];
assign w281 = ~in10[2];
assign w282 = ~in10[2];
assign w283 = ~in10[2];
assign w284 = ~in10[3];
assign w285 = ~in10[3];
assign w286 = ~in10[3];
assign w287 = ~in10[3];
assign w288 = ~in10[3];
assign w289 = ~in10[3];
assign w290 = in1[10] & in10[4];
assign w291 = ~in10[4];
assign w292 = ~in10[4];
assign w293 = ~in10[4];
assign w294 = ~in10[4];
assign w295 = ~in10[4];
assign w296 = ~in10[4];
assign w297 = ~in11[1];
assign w298 = w11 ~^ in1[2];
assign w299 = in1[0] | w12;
assign w300 = w11 | w15;
assign w301 = w18 ~^ in1[4];
assign w302 = w18 | w21;
assign w303 = w24 ~^ in1[6];
assign w304 = w24 | w27;
assign w305 = w30 ~^ in1[8];
assign w306 = w30 | w33;
assign w307 = w36 ~^ in1[10];
assign w308 = w36 | w39;
assign w309 = ~w44;
assign w310 = ~w44;
assign w311 = ~w44;
assign w312 = ~w44;
assign w313 = ~w44;
assign w314 = ~w44;
assign w315 = ~w44;
assign w316 = ~w44;
assign w317 = w3 | w50;
assign w318 = w4 | w56;
assign w319 = w2 | w62;
assign w320 = w1 | w68;
assign w321 = w6 | w74;
assign w322 = w1 | w80;
assign w323 = w2 | w86;
assign w324 = w44 ~| w88;
assign w325 = w5 | w93;
assign w326 = w44 | w95;
assign w327 = w3 | w100;
assign w328 = w7 | w105;
assign w329 = w7 | w112;
assign w330 = w8 | w118;
assign w331 = w5 | w123;
assign w332 = w4 | w130;
assign w333 = w6 | w136;
assign w334 = w8 | w142;
assign w335 = w1 | w148;
assign w336 = w44 ~| w150;
assign w337 = w167 | w170;
assign w338 = w171 | w174;
assign w339 = w175 | w178;
assign w340 = w183 | w186;
assign w341 = ~w187;
assign w342 = w205 | in4;
assign w343 = w203 & w205;
assign w344 = w204 & w206;
assign w345 = w214 ~| in9[31];
assign w346 = w215 ~| in9[0];
assign w347 = w217 ~| in9[17];
assign w348 = w218 ~| in9[25];
assign w349 = w218 ~| in9[27];
assign w350 = w219 ~| in9[21];
assign w351 = w219 ~| in9[23];
assign w352 = w221 ~| in9[24];
assign w353 = w238 ~| in9[19];
assign w354 = w239 ~| in9[18];
assign w355 = w241 ~| in9[22];
assign w356 = w243 ~| in9[26];
assign w357 = w243 ~| in9[28];
assign w358 = w244 ~| in9[20];
assign w359 = w245 ~| in9[29];
assign w360 = w245 ~| in9[30];
assign w361 = w217 ~| w263;
assign w362 = w37 | w264;
assign w363 = w22 | w264;
assign w364 = w28 | w264;
assign w365 = w34 | w265;
assign w366 = w16 | w265;
assign w367 = w31 | w266;
assign w368 = w25 | w266;
assign w369 = w40 | w267;
assign w370 = w13 | w268;
assign w371 = w19 | w268;
assign w372 = w43 | w269;
assign w373 = w37 | w270;
assign w374 = w28 | w270;
assign w375 = w16 | w270;
assign w376 = w34 | w271;
assign w377 = w31 | w271;
assign w378 = w0 | w271;
assign w379 = w43 | w272;
assign w380 = w25 | w272;
assign w381 = w9 | w273;
assign w382 = w19 | w273;
assign w383 = w40 | w274;
assign w384 = w22 | w274;
assign w385 = w13 | w275;
assign w386 = in9[8] ~| w276;
assign w387 = ~w276;
assign w388 = in9[9] ~| w277;
assign w389 = ~w277;
assign w390 = in9[7] ~| w278;
assign w391 = ~w278;
assign w392 = w34 | w279;
assign w393 = w9 | w279;
assign w394 = w0 | w280;
assign w395 = w31 | w280;
assign w396 = w43 | w280;
assign w397 = w19 | w281;
assign w398 = w16 | w281;
assign w399 = w40 | w282;
assign w400 = w13 | w282;
assign w401 = w37 | w283;
assign w402 = w0 | w284;
assign w403 = w22 | w284;
assign w404 = w28 | w284;
assign w405 = w40 | w285;
assign w406 = w43 | w285;
assign w407 = w9 | w285;
assign w408 = w19 | w286;
assign w409 = w13 | w286;
assign w410 = w37 | w287;
assign w411 = w34 | w287;
assign w412 = w25 | w288;
assign w413 = w31 | w288;
assign w414 = w16 | w289;
assign w415 = in9[14] ~| w290;
assign w416 = ~w290;
assign w417 = w28 | w291;
assign w418 = w43 | w291;
assign w419 = w31 | w291;
assign w420 = w34 | w292;
assign w421 = w19 | w292;
assign w422 = w0 | w292;
assign w423 = w40 | w293;
assign w424 = w16 | w293;
assign w425 = w9 | w294;
assign w426 = w25 | w295;
assign w427 = w13 | w295;
assign w428 = w22 | w296;
assign w429 = ~w298;
assign w430 = ~w298;
assign w431 = ~w298;
assign w432 = in1[3] & w298;
assign w433 = w17 | w298;
assign w434 = ~w298;
assign w435 = ~w298;
assign w436 = ~w298;
assign w437 = ~w298;
assign w438 = ~w298;
assign w439 = ~w298;
assign w440 = w148 ~| w299;
assign w441 = w136 | w299;
assign w442 = w142 | w299;
assign w443 = w130 | w299;
assign w444 = w112 | w299;
assign w445 = w74 | w299;
assign w446 = w118 | w299;
assign w447 = w11 ~| w299;
assign w448 = w62 | w299;
assign w449 = w50 | w299;
assign w450 = w123 | w299;
assign w451 = w100 | w299;
assign w452 = w80 | w299;
assign w453 = w68 | w299;
assign w454 = w56 | w299;
assign w455 = w105 | w299;
assign w456 = w93 | w299;
assign w457 = in2[0] | w299;
assign w458 = w86 | w299;
assign w459 = ~w301;
assign w460 = ~w301;
assign w461 = ~w301;
assign w462 = in1[5] & w301;
assign w463 = w23 | w301;
assign w464 = ~w301;
assign w465 = ~w301;
assign w466 = ~w301;
assign w467 = ~w301;
assign w468 = ~w301;
assign w469 = ~w301;
assign w470 = ~w303;
assign w471 = ~w303;
assign w472 = ~w303;
assign w473 = in1[7] & w303;
assign w474 = w29 | w303;
assign w475 = ~w303;
assign w476 = ~w303;
assign w477 = ~w303;
assign w478 = ~w303;
assign w479 = ~w303;
assign w480 = ~w303;
assign w481 = ~w305;
assign w482 = ~w305;
assign w483 = ~w305;
assign w484 = in1[9] & w305;
assign w485 = w35 | w305;
assign w486 = ~w305;
assign w487 = ~w305;
assign w488 = ~w305;
assign w489 = ~w305;
assign w490 = ~w305;
assign w491 = ~w305;
assign w492 = ~w307;
assign w493 = ~w307;
assign w494 = ~w307;
assign w495 = in1[11] & w307;
assign w496 = w41 | w307;
assign w497 = ~w307;
assign w498 = ~w307;
assign w499 = ~w307;
assign w500 = ~w307;
assign w501 = ~w307;
assign w502 = ~w307;
assign w503 = in2[2] & w309;
assign w504 = w45 | w309;
assign w505 = in2[11] & w310;
assign w506 = in2[1] & w310;
assign w507 = in2[5] & w311;
assign w508 = in2[3] & w312;
assign w509 = in2[4] & w312;
assign w510 = in2[14] & w313;
assign w511 = in2[10] & w313;
assign w512 = in2[16] & w314;
assign w513 = in2[12] & w314;
assign w514 = in2[13] & w315;
assign w515 = in2[15] & w315;
assign w516 = in2[6] & w316;
assign w517 = in2[9] & w316;
assign w518 = ~w342;
assign w519 = ~w342;
assign w520 = ~w342;
assign w521 = ~w342;
assign w522 = ~w342;
assign w523 = ~w342;
assign w524 = ~w342;
assign w525 = ~w342;
assign w526 = ~w342;
assign w527 = ~w342;
assign w528 = ~w342;
assign w529 = ~w342;
assign w530 = ~w342;
assign w531 = ~w342;
assign w532 = ~w342;
assign w533 = ~w342;
assign w534 = ~w343;
assign w535 = ~w343;
assign w536 = ~w343;
assign w537 = ~w343;
assign w538 = ~w343;
assign w539 = ~w343;
assign w540 = ~w343;
assign w541 = ~w343;
assign w542 = ~w343;
assign w543 = ~w343;
assign w544 = ~w343;
assign w545 = ~w343;
assign w546 = ~w343;
assign w547 = ~w343;
assign w548 = ~w343;
assign w549 = ~w343;
assign w550 = ~w344;
assign w551 = ~w344;
assign w552 = ~w344;
assign w553 = ~w344;
assign w554 = ~w344;
assign w555 = ~w344;
assign w556 = ~w344;
assign w557 = ~w344;
assign w558 = ~w344;
assign w559 = ~w344;
assign w560 = ~w344;
assign w561 = ~w344;
assign w562 = w362 ~^ in9[10];
assign w563 = w363 ~^ in9[5];
assign w564 = w364 ~^ in9[7];
assign w565 = w365 ~^ in9[9];
assign w566 = w366 ~^ in9[3];
assign w567 = ~w366;
assign w568 = w367 ~^ in9[8];
assign w569 = w368 ~^ in9[6];
assign w570 = w369 ~^ in9[11];
assign w571 = w370 ~^ in9[2];
assign w572 = w189 | w370;
assign w573 = w371 ~^ in9[4];
assign w574 = w190 | w371;
assign w575 = w372 ~^ in9[12];
assign w576 = w378 ~^ in9[1];
assign w577 = ~w378;
assign w578 = w379 ~^ in9[13];
assign w579 = w199 | w379;
assign w580 = ~w381;
assign w581 = w367 | w386;
assign w582 = w194 | w387;
assign w583 = w365 | w388;
assign w584 = w195 | w389;
assign w585 = w364 | w390;
assign w586 = w193 | w391;
assign w587 = w197 | w392;
assign w588 = ~w392;
assign w589 = w381 ~^ w394;
assign w590 = w381 ~| w394;
assign w591 = ~w394;
assign w592 = w196 | w395;
assign w593 = ~w395;
assign w594 = w396 ~^ in9[14];
assign w595 = w192 | w397;
assign w596 = ~w397;
assign w597 = w191 | w398;
assign w598 = ~w398;
assign w599 = w198 & w401;
assign w600 = w198 ~| w401;
assign w601 = w393 ~^ w402;
assign w602 = w393 & w402;
assign w603 = w393 | w402;
assign w604 = w374 ~^ w403;
assign w605 = w376 ~^ w404;
assign w606 = w406 ~^ in9[15];
assign w607 = w400 ~^ w407;
assign w608 = w400 & w407;
assign w609 = w400 | w407;
assign w610 = w380 ~^ w408;
assign w611 = w382 ~^ w409;
assign w612 = w383 ~^ w411;
assign w613 = w377 ~^ w412;
assign w614 = w373 ~^ w413;
assign w615 = w384 ~^ w414;
assign w616 = w396 | w415;
assign w617 = w200 | w416;
assign w618 = w413 & w417;
assign w619 = w413 | w417;
assign w620 = w418 ~^ in9[16];
assign w621 = w202 ~| w418;
assign w622 = w202 & w418;
assign w623 = w411 & w419;
assign w624 = w411 | w419;
assign w625 = w410 ~^ w420;
assign w626 = w410 | w420;
assign w627 = w410 & w420;
assign w628 = w403 | w421;
assign w629 = w403 & w421;
assign w630 = ~w422;
assign w631 = w201 | w423;
assign w632 = ~w423;
assign w633 = w408 | w424;
assign w634 = w408 & w424;
assign w635 = w409 & w425;
assign w636 = w409 | w425;
assign w637 = w404 | w426;
assign w638 = w404 & w426;
assign w639 = w414 | w427;
assign w640 = w414 & w427;
assign w641 = w412 & w428;
assign w642 = w412 | w428;
assign w643 = w85 | w429;
assign w644 = w53 | w429;
assign w645 = w117 | w430;
assign w646 = w128 | w430;
assign w647 = w97 | w431;
assign w648 = w146 | w431;
assign w649 = w91 | w431;
assign w650 = ~w432;
assign w651 = w135 | w433;
assign w652 = w47 | w433;
assign w653 = w66 | w433;
assign w654 = w108 | w433;
assign w655 = w146 | w433;
assign w656 = w103 | w433;
assign w657 = w18 ~| w433;
assign w658 = w117 | w433;
assign w659 = w128 | w433;
assign w660 = w79 | w433;
assign w661 = w85 | w433;
assign w662 = w91 | w433;
assign w663 = w53 | w433;
assign w664 = w122 | w433;
assign w665 = w97 | w433;
assign w666 = w73 | w433;
assign w667 = w140 | w433;
assign w668 = w60 | w433;
assign w669 = w60 | w434;
assign w670 = w47 | w434;
assign w671 = w135 | w435;
assign w672 = w140 | w436;
assign w673 = w79 | w436;
assign w674 = w66 | w437;
assign w675 = w103 | w438;
assign w676 = w73 | w438;
assign w677 = w122 | w439;
assign w678 = w108 | w439;
assign w679 = w10 | w440;
assign w680 = w334 & w441;
assign w681 = w335 & w442;
assign w682 = w333 & w443;
assign w683 = w330 & w444;
assign w684 = w322 & w445;
assign w685 = w331 & w446;
assign w686 = w10 | w447;
assign w687 = w320 & w448;
assign w688 = w318 & w449;
assign w689 = w332 & w450;
assign w690 = w328 & w451;
assign w691 = w323 & w452;
assign w692 = w321 & w453;
assign w693 = w319 & w454;
assign w694 = w329 & w455;
assign w695 = w327 & w456;
assign w696 = w317 & w457;
assign w697 = w325 & w458;
assign w698 = w70 | w459;
assign w699 = w49 | w459;
assign w700 = w145 | w460;
assign w701 = w127 | w460;
assign w702 = w111 | w461;
assign w703 = w99 | w461;
assign w704 = w124 | w461;
assign w705 = ~w462;
assign w706 = w90 | w463;
assign w707 = w133 | w463;
assign w708 = w127 | w463;
assign w709 = w70 | w463;
assign w710 = w102 | w463;
assign w711 = w49 | w463;
assign w712 = w124 | w463;
assign w713 = w24 ~| w463;
assign w714 = w84 | w463;
assign w715 = w114 | w463;
assign w716 = w99 | w463;
assign w717 = w111 | w463;
assign w718 = w138 | w463;
assign w719 = w145 | w463;
assign w720 = w59 | w463;
assign w721 = w52 | w463;
assign w722 = w64 | w463;
assign w723 = w78 | w463;
assign w724 = w90 | w464;
assign w725 = w114 | w464;
assign w726 = w52 | w465;
assign w727 = w133 | w466;
assign w728 = w102 | w466;
assign w729 = w84 | w467;
assign w730 = w138 | w468;
assign w731 = w78 | w468;
assign w732 = w59 | w469;
assign w733 = w64 | w469;
assign w734 = w46 | w470;
assign w735 = w147 | w470;
assign w736 = w61 | w471;
assign w737 = w77 | w471;
assign w738 = w120 | w472;
assign w739 = w92 | w472;
assign w740 = w55 | w472;
assign w741 = ~w473;
assign w742 = w65 | w474;
assign w743 = w134 | w474;
assign w744 = w55 | w474;
assign w745 = w147 | w474;
assign w746 = w96 | w474;
assign w747 = w120 | w474;
assign w748 = w116 | w474;
assign w749 = w30 ~| w474;
assign w750 = w83 | w474;
assign w751 = w110 | w474;
assign w752 = w46 | w474;
assign w753 = w129 | w474;
assign w754 = w106 | w474;
assign w755 = w77 | w474;
assign w756 = w72 | w474;
assign w757 = w61 | w474;
assign w758 = w139 | w474;
assign w759 = w92 | w474;
assign w760 = w72 | w475;
assign w761 = w65 | w475;
assign w762 = w106 | w476;
assign w763 = w110 | w477;
assign w764 = w83 | w477;
assign w765 = w139 | w478;
assign w766 = w134 | w479;
assign w767 = w116 | w479;
assign w768 = w129 | w480;
assign w769 = w96 | w480;
assign w770 = w115 | w481;
assign w771 = w141 | w481;
assign w772 = w89 | w482;
assign w773 = w82 | w482;
assign w774 = w71 | w483;
assign w775 = w121 | w483;
assign w776 = w58 | w483;
assign w777 = ~w484;
assign w778 = w54 | w485;
assign w779 = w48 | w485;
assign w780 = w144 | w485;
assign w781 = w121 | w485;
assign w782 = w82 | w485;
assign w783 = w132 | w485;
assign w784 = w36 ~| w485;
assign w785 = w109 | w485;
assign w786 = w76 | w485;
assign w787 = w104 | w485;
assign w788 = w115 | w485;
assign w789 = w71 | w485;
assign w790 = w89 | w485;
assign w791 = w126 | w485;
assign w792 = w58 | w485;
assign w793 = w98 | w485;
assign w794 = w67 | w485;
assign w795 = w141 | w485;
assign w796 = w132 | w486;
assign w797 = w109 | w486;
assign w798 = w104 | w487;
assign w799 = w54 | w488;
assign w800 = w144 | w488;
assign w801 = w76 | w489;
assign w802 = w48 | w490;
assign w803 = w98 | w490;
assign w804 = w126 | w491;
assign w805 = w67 | w491;
assign w806 = w137 | w492;
assign w807 = w113 | w492;
assign w808 = w107 | w493;
assign w809 = w119 | w493;
assign w810 = w57 | w494;
assign w811 = w149 | w494;
assign w812 = w87 | w494;
assign w813 = ~w495;
assign w814 = w125 | w496;
assign w815 = w69 | w496;
assign w816 = w101 | w496;
assign w817 = w131 | w496;
assign w818 = w137 | w496;
assign w819 = w81 | w496;
assign w820 = w63 | w496;
assign w821 = w42 ~| w496;
assign w822 = w107 | w496;
assign w823 = w149 | w496;
assign w824 = w143 | w496;
assign w825 = w75 | w496;
assign w826 = w57 | w496;
assign w827 = w119 | w496;
assign w828 = w94 | w496;
assign w829 = w87 | w496;
assign w830 = w51 | w496;
assign w831 = w113 | w496;
assign w832 = w69 | w497;
assign w833 = w131 | w497;
assign w834 = w125 | w498;
assign w835 = w75 | w499;
assign w836 = w101 | w499;
assign w837 = w143 | w500;
assign w838 = w63 | w501;
assign w839 = w94 | w501;
assign w840 = w51 | w502;
assign w841 = w81 | w502;
assign w842 = ~w504;
assign w843 = ~w504;
assign w844 = ~w504;
assign w845 = ~w504;
assign w846 = w88 | w504;
assign w847 = w150 | w504;
assign w848 = ~w504;
assign w849 = ~w504;
assign w850 = ~w504;
assign w851 = w254 | w534;
assign w852 = w253 | w534;
assign w853 = w249 | w535;
assign w854 = w227 | w535;
assign w855 = w230 | w536;
assign w856 = w256 | w536;
assign w857 = w235 | w537;
assign w858 = w258 | w537;
assign w859 = w237 | w538;
assign w860 = w261 | w538;
assign w861 = w233 | w539;
assign w862 = w246 | w539;
assign w863 = w232 | w540;
assign w864 = w223 | w540;
assign w865 = w228 | w541;
assign w866 = w226 | w541;
assign w867 = w225 | w542;
assign w868 = w250 | w542;
assign w869 = w259 | w543;
assign w870 = w248 | w543;
assign w871 = w222 | w544;
assign w872 = w231 | w544;
assign w873 = w229 | w545;
assign w874 = w251 | w545;
assign w875 = w224 | w546;
assign w876 = w255 | w546;
assign w877 = w234 | w547;
assign w878 = w252 | w547;
assign w879 = w257 | w548;
assign w880 = w236 | w548;
assign w881 = w260 | w549;
assign w882 = w247 | w549;
assign w883 = w209 ~| w550;
assign w884 = w209 ~| w551;
assign w885 = w211 ~| w552;
assign w886 = w211 ~| w553;
assign w887 = w211 ~| w554;
assign w888 = w210 ~| w554;
assign w889 = w210 ~| w555;
assign w890 = w211 ~| w555;
assign w891 = w207 ~| w556;
assign w892 = w208 ~| w556;
assign w893 = w207 ~| w557;
assign w894 = w208 ~| w557;
assign w895 = w207 ~| w558;
assign w896 = w208 ~| w559;
assign w897 = w213 ~| w560;
assign w898 = w212 ~| w560;
assign w899 = w212 ~| w561;
assign w900 = w213 ~| w561;
assign w901 = w395 ~^ w562;
assign w902 = w398 ~^ w563;
assign w903 = w391 ~^ w564;
assign w904 = w389 ~^ w565;
assign w905 = ~w566;
assign w906 = in9[3] & w567;
assign w907 = w387 ~^ w568;
assign w908 = w397 ~^ w569;
assign w909 = w392 ~^ w570;
assign w910 = w566 ~^ w572;
assign w911 = w422 ~^ w573;
assign w912 = w401 ~^ w575;
assign w913 = in9[1] & w577;
assign w914 = ~w578;
assign w915 = w405 ~^ w579;
assign w916 = w405 | w579;
assign w917 = w405 & w579;
assign w918 = w581 & w582;
assign w919 = w583 & w584;
assign w920 = w585 & w586;
assign w921 = in9[11] ~| w588;
assign w922 = w571 ~^ w589;
assign w923 = w580 | w591;
assign w924 = in9[10] ~| w593;
assign w925 = w416 ~^ w594;
assign w926 = in9[6] ~| w596;
assign w927 = in9[5] ~| w598;
assign w928 = w372 ~| w599;
assign w929 = w385 ~^ w601;
assign w930 = w385 | w602;
assign w931 = w421 ~^ w604;
assign w932 = w426 ~^ w605;
assign w933 = w423 ~^ w606;
assign w934 = w375 ~^ w607;
assign w935 = w375 | w608;
assign w936 = w424 ~^ w610;
assign w937 = w425 ~^ w611;
assign w938 = w419 ~^ w612;
assign w939 = w428 ~^ w613;
assign w940 = w417 ~^ w614;
assign w941 = w427 ~^ w615;
assign w942 = w616 & w617;
assign w943 = w373 | w618;
assign w944 = w383 | w623;
assign w945 = w399 ~^ w625;
assign w946 = w399 | w627;
assign w947 = w374 | w629;
assign w948 = in9[15] ~| w632;
assign w949 = w380 | w634;
assign w950 = w382 | w635;
assign w951 = w376 | w638;
assign w952 = w384 | w640;
assign w953 = w377 | w641;
assign w954 = w644 & w652;
assign w955 = w645 & w654;
assign w956 = w650 & w655;
assign w957 = w432 | w657;
assign w958 = w643 & w660;
assign w959 = w649 & w661;
assign w960 = w647 & w662;
assign w961 = w646 & w664;
assign w962 = w648 & w667;
assign w963 = w663 & w669;
assign w964 = w659 & w671;
assign w965 = w651 & w672;
assign w966 = w666 & w673;
assign w967 = w668 & w674;
assign w968 = w665 & w675;
assign w969 = w653 & w676;
assign w970 = w658 & w677;
assign w971 = w656 & w678;
assign w972 = w679 ~^ in3[18];
assign w973 = ~w679;
assign w974 = w680 ~^ in3[16];
assign w975 = ~w680;
assign w976 = w681 ~^ in3[17];
assign w977 = w164 | w681;
assign w978 = w682 ~^ in3[15];
assign w979 = ~w682;
assign w980 = w685 ~^ in3[13];
assign w981 = ~w687;
assign w982 = w689 ~^ in3[14];
assign w983 = ~w689;
assign w984 = ~w697;
assign w985 = w703 & w706;
assign w986 = w702 & w710;
assign w987 = w701 & w712;
assign w988 = w462 | w713;
assign w989 = w704 & w715;
assign w990 = w700 & w718;
assign w991 = w705 & w719;
assign w992 = w698 & w722;
assign w993 = w714 & w724;
assign w994 = w717 & w725;
assign w995 = w711 & w726;
assign w996 = w708 & w727;
assign w997 = w716 & w728;
assign w998 = w723 & w729;
assign w999 = w707 & w730;
assign w1000 = w709 & w731;
assign w1001 = w721 & w732;
assign w1002 = w720 & w733;
assign w1003 = w736 & w744;
assign w1004 = w741 & w745;
assign w1005 = w738 & w748;
assign w1006 = w473 | w749;
assign w1007 = w739 & w750;
assign w1008 = w740 & w752;
assign w1009 = w737 & w756;
assign w1010 = w735 & w758;
assign w1011 = w742 & w760;
assign w1012 = w757 & w761;
assign w1013 = w746 & w762;
assign w1014 = w754 & w763;
assign w1015 = w755 & w764;
assign w1016 = w743 & w765;
assign w1017 = w753 & w766;
assign w1018 = w751 & w767;
assign w1019 = w747 & w768;
assign w1020 = w759 & w769;
assign w1021 = w776 & w778;
assign w1022 = w777 & w780;
assign w1023 = w772 & w782;
assign w1024 = w771 & w783;
assign w1025 = w484 | w784;
assign w1026 = w770 & w785;
assign w1027 = w773 & w786;
assign w1028 = w775 & w788;
assign w1029 = w774 & w794;
assign w1030 = w791 & w796;
assign w1031 = w787 & w797;
assign w1032 = w793 & w798;
assign w1033 = w779 & w799;
assign w1034 = w795 & w800;
assign w1035 = w789 & w801;
assign w1036 = w790 & w803;
assign w1037 = w781 & w804;
assign w1038 = w792 & w805;
assign w1039 = w808 & w816;
assign w1040 = w806 & w817;
assign w1041 = w812 & w819;
assign w1042 = w495 | w821;
assign w1043 = w807 & w822;
assign w1044 = w813 & w823;
assign w1045 = w811 & w824;
assign w1046 = w810 & w830;
assign w1047 = w809 & w831;
assign w1048 = w820 & w832;
assign w1049 = w814 & w833;
assign w1050 = w827 & w834;
assign w1051 = w815 & w835;
assign w1052 = w828 & w836;
assign w1053 = w818 & w837;
assign w1054 = w826 & w838;
assign w1055 = w829 & w839;
assign w1056 = w825 & w841;
assign w1057 = in2[12] & w842;
assign w1058 = in2[4] & w842;
assign w1059 = in2[2] & w843;
assign w1060 = in2[15] & w843;
assign w1061 = in2[11] & w844;
assign w1062 = in2[16] & w844;
assign w1063 = in2[5] & w845;
assign w1064 = in2[10] & w845;
assign w1065 = w326 & w846;
assign w1066 = w847 ~^ in3[30];
assign w1067 = in3[30] & w847;
assign w1068 = in3[30] | w847;
assign w1069 = in2[6] & w848;
assign w1070 = in2[14] & w848;
assign w1071 = in2[3] & w848;
assign w1072 = in2[13] & w849;
assign w1073 = in2[9] & w849;
assign w1074 = in2[1] & w850;
assign w1075 = in2[8] & w850;
assign w1076 = w345 ~| w852;
assign w1077 = w361 ~| w855;
assign w1078 = w346 ~| w857;
assign w1079 = w349 ~| w858;
assign w1080 = w357 ~| w859;
assign w1081 = w355 ~| w860;
assign w1082 = w359 ~| w861;
assign w1083 = w356 ~| w862;
assign w1084 = w350 ~| w863;
assign w1085 = w354 ~| w865;
assign w1086 = w348 ~| w867;
assign w1087 = w360 ~| w868;
assign w1088 = w352 ~| w872;
assign w1089 = w353 ~| w878;
assign w1090 = w358 ~| w879;
assign w1091 = w347 ~| w881;
assign w1092 = w351 ~| w882;
assign w1093 = w262 & w890;
assign w1094 = w576 & w899;
assign w1095 = ~w901;
assign w1096 = ~w902;
assign w1097 = ~w903;
assign w1098 = ~w904;
assign w1099 = w572 ~| w905;
assign w1100 = w572 & w905;
assign w1101 = w630 | w906;
assign w1102 = ~w906;
assign w1103 = ~w907;
assign w1104 = ~w908;
assign w1105 = ~w909;
assign w1106 = ~w912;
assign w1107 = w214 ~| w913;
assign w1108 = w369 | w921;
assign w1109 = w883 & w922;
assign w1110 = w571 & w923;
assign w1111 = w362 | w924;
assign w1112 = ~w925;
assign w1113 = w368 | w926;
assign w1114 = w363 | w927;
assign w1115 = w600 | w928;
assign w1116 = w910 ~^ w929;
assign w1117 = w603 & w930;
assign w1118 = ~w933;
assign w1119 = ~w934;
assign w1120 = w609 & w935;
assign w1121 = ~w937;
assign w1122 = w933 ~^ w942;
assign w1123 = w619 & w943;
assign w1124 = w624 & w944;
assign w1125 = w626 & w946;
assign w1126 = w628 & w947;
assign w1127 = w406 | w948;
assign w1128 = w633 & w949;
assign w1129 = w636 & w950;
assign w1130 = w637 & w951;
assign w1131 = w639 & w952;
assign w1132 = w642 & w953;
assign w1133 = w687 ~^ w954;
assign w1134 = w687 ~| w954;
assign w1135 = ~w954;
assign w1136 = in3[20] & w956;
assign w1137 = in3[20] | w956;
assign w1138 = w168 ~^ w957;
assign w1139 = w169 | w957;
assign w1140 = w691 ~^ w969;
assign w1141 = w691 & w969;
assign w1142 = w691 ~| w969;
assign w1143 = w165 | w973;
assign w1144 = ~w974;
assign w1145 = in3[16] & w975;
assign w1146 = ~w976;
assign w1147 = w972 ~^ w977;
assign w1148 = w972 | w977;
assign w1149 = w972 & w977;
assign w1150 = ~w978;
assign w1151 = in3[15] & w979;
assign w1152 = ~w982;
assign w1153 = in3[14] & w983;
assign w1154 = ~w986;
assign w1155 = ~w987;
assign w1156 = w172 ~^ w988;
assign w1157 = w173 | w988;
assign w1158 = ~w994;
assign w1159 = w996 ~^ in3[19];
assign w1160 = w166 & w996;
assign w1161 = ~w997;
assign w1162 = w992 ~^ w1003;
assign w1163 = ~w1005;
assign w1164 = w176 ~^ w1006;
assign w1165 = w177 | w1006;
assign w1166 = w955 ~^ w1007;
assign w1167 = w955 & w1007;
assign w1168 = w955 | w1007;
assign w1169 = w966 ~^ w1008;
assign w1170 = w960 ~^ w1011;
assign w1171 = w960 | w1011;
assign w1172 = w960 & w1011;
assign w1173 = w985 ~^ w1015;
assign w1174 = w985 | w1015;
assign w1175 = w985 & w1015;
assign w1176 = ~w1016;
assign w1177 = w961 ~^ w1023;
assign w1178 = w961 | w1023;
assign w1179 = w961 & w1023;
assign w1180 = w1019 ~^ w1026;
assign w1181 = w970 ~^ w1027;
assign w1182 = w970 | w1027;
assign w1183 = w970 & w1027;
assign w1184 = w1017 ~^ w1028;
assign w1185 = w1017 & w1028;
assign w1186 = w1017 | w1028;
assign w1187 = ~w1030;
assign w1188 = w962 ~^ w1031;
assign w1189 = w965 ~^ w1032;
assign w1190 = w690 ~^ w1033;
assign w1191 = w690 | w1033;
assign w1192 = w690 & w1033;
assign w1193 = w964 ~^ w1036;
assign w1194 = w1037 ~^ in3[22];
assign w1195 = w968 ~^ w1038;
assign w1196 = w968 | w1038;
assign w1197 = w968 & w1038;
assign w1198 = w1026 & w1039;
assign w1199 = w1026 | w1039;
assign w1200 = ~w1040;
assign w1201 = w964 | w1041;
assign w1202 = w964 & w1041;
assign w1203 = w184 ~^ w1042;
assign w1204 = w185 | w1042;
assign w1205 = ~w1043;
assign w1206 = w1025 ~^ w1045;
assign w1207 = w1025 & w1045;
assign w1208 = w1025 | w1045;
assign w1209 = in3[22] | w1047;
assign w1210 = in3[22] & w1047;
assign w1211 = w982 ~^ w1048;
assign w1212 = ~w1048;
assign w1213 = w1024 ~^ w1049;
assign w1214 = w1024 | w1049;
assign w1215 = w1024 & w1049;
assign w1216 = w1030 ~^ w1050;
assign w1217 = w1031 & w1052;
assign w1218 = w1031 | w1052;
assign w1219 = w1029 ~^ w1054;
assign w1220 = w1029 | w1054;
assign w1221 = w1029 & w1054;
assign w1222 = w965 | w1055;
assign w1223 = w965 & w1055;
assign w1224 = w514 | w1057;
assign w1225 = w507 | w1058;
assign w1226 = w508 | w1059;
assign w1227 = w512 | w1060;
assign w1228 = w513 | w1061;
assign w1229 = w336 | w1062;
assign w1230 = w516 | w1063;
assign w1231 = w505 | w1064;
assign w1232 = w1065 ^ in3[20];
assign w1233 = w324 | w1069;
assign w1234 = w515 | w1070;
assign w1235 = w509 | w1071;
assign w1236 = w510 | w1072;
assign w1237 = w511 | w1073;
assign w1238 = w503 | w1074;
assign w1239 = w517 | w1075;
assign w1240 = w1094 ~^ in11[1];
assign w1241 = ~w1094;
assign w1242 = w929 ~| w1100;
assign w1243 = w573 & w1101;
assign w1244 = w911 ~^ w1102;
assign w1245 = w422 ~| w1102;
assign w1246 = w873 ~| w1107;
assign w1247 = w587 & w1108;
assign w1248 = w1109;
assign w1249 = w590 | w1110;
assign w1250 = w592 & w1111;
assign w1251 = w595 & w1113;
assign w1252 = w597 & w1114;
assign w1253 = w578 ~| w1115;
assign w1254 = ~w1115;
assign w1255 = w1116;
assign w1256 = w934 ~^ w1117;
assign w1257 = w934 ~| w1117;
assign w1258 = ~w1117;
assign w1259 = w942 & w1118;
assign w1260 = w942 ~| w1118;
assign w1261 = w574 ~^ w1120;
assign w1262 = w574 | w1120;
assign w1263 = w574 & w1120;
assign w1264 = w915 ~^ w1125;
assign w1265 = w917 | w1125;
assign w1266 = w1098 | w1126;
assign w1267 = w918 ~^ w1126;
assign w1268 = ~w1126;
assign w1269 = w631 & w1127;
assign w1270 = w1103 | w1128;
assign w1271 = w920 ~^ w1128;
assign w1272 = ~w1128;
assign w1273 = w1097 | w1131;
assign w1274 = ~w1131;
assign w1275 = w1095 | w1132;
assign w1276 = w919 ~^ w1132;
assign w1277 = ~w1132;
assign w1278 = w981 | w1135;
assign w1279 = w1065 | w1136;
assign w1280 = w337 & w1139;
assign w1281 = w976 ~| w1145;
assign w1282 = ~w1145;
assign w1283 = w974 ~| w1151;
assign w1284 = ~w1151;
assign w1285 = w1048 ~| w1152;
assign w1286 = ~w1153;
assign w1287 = ~w1156;
assign w1288 = w338 & w1157;
assign w1289 = w1143 ~^ w1159;
assign w1290 = w1143 & w1159;
assign w1291 = w1143 | w1159;
assign w1292 = w999 ~^ w1160;
assign w1293 = w999 | w1160;
assign w1294 = w999 & w1160;
assign w1295 = ~w1164;
assign w1296 = w339 & w1165;
assign w1297 = w1035 ~^ w1166;
assign w1298 = w1035 | w1167;
assign w1299 = w1021 ~^ w1170;
assign w1300 = w1021 | w1172;
assign w1301 = w971 ~^ w1173;
assign w1302 = w971 | w1175;
assign w1303 = w1056 ~^ w1177;
assign w1304 = w1056 | w1179;
assign w1305 = w1039 ~^ w1180;
assign w1306 = w1051 ~^ w1181;
assign w1307 = w1051 | w1183;
assign w1308 = w990 ~^ w1184;
assign w1309 = w990 | w1185;
assign w1310 = w1052 ~^ w1188;
assign w1311 = w1055 ~^ w1189;
assign w1312 = w1041 ~^ w1193;
assign w1313 = w1047 ~^ w1194;
assign w1314 = w1046 ~^ w1195;
assign w1315 = w1046 | w1197;
assign w1316 = w1019 | w1198;
assign w1317 = w1036 | w1202;
assign w1318 = ~w1203;
assign w1319 = w340 & w1204;
assign w1320 = w1037 | w1210;
assign w1321 = w982 | w1212;
assign w1322 = w962 | w1217;
assign w1323 = w1032 | w1223;
assign w1324 = w1040 ~^ w1224;
assign w1325 = w1200 ~| w1224;
assign w1326 = ~w1224;
assign w1327 = w989 ~^ w1225;
assign w1328 = ~w1225;
assign w1329 = w986 ~^ w1226;
assign w1330 = w1154 ~| w1226;
assign w1331 = ~w1226;
assign w1332 = w1227 ~^ in3[28];
assign w1333 = w183 ~| w1227;
assign w1334 = ~w1227;
assign w1335 = w1228 ~^ in3[24];
assign w1336 = w175 ~| w1228;
assign w1337 = ~w1228;
assign w1338 = w1203 ~^ w1229;
assign w1339 = ~w1229;
assign w1340 = w987 ~^ w1230;
assign w1341 = w1155 ~| w1230;
assign w1342 = ~w1230;
assign w1343 = w1216 ~^ w1231;
assign w1344 = w1187 ~| w1231;
assign w1345 = ~w1231;
assign w1346 = w956 ~^ w1232;
assign w1347 = w686 ~^ w1233;
assign w1348 = w1163 ~| w1233;
assign w1349 = ~w1233;
assign w1350 = w180 ~^ w1234;
assign w1351 = w182 & w1234;
assign w1352 = w994 ~^ w1235;
assign w1353 = w1158 ~| w1235;
assign w1354 = ~w1235;
assign w1355 = w1236 ~^ in3[26];
assign w1356 = w179 ~| w1236;
assign w1357 = ~w1236;
assign w1358 = w991 ~^ w1237;
assign w1359 = w1176 ~| w1237;
assign w1360 = ~w1237;
assign w1361 = w997 ~^ w1238;
assign w1362 = w1161 & w1238;
assign w1363 = w1043 ~^ w1239;
assign w1364 = w1205 ~| w1239;
assign w1365 = ~w1239;
assign w1366 = ~w1240;
assign w1367 = w297 | w1241;
assign w1368 = w1099 | w1242;
assign w1369 = w1243 | w1245;
assign w1370 = w1123 ~^ w1247;
assign w1371 = w1123 & w1247;
assign w1372 = w1123 | w1247;
assign w1373 = w1248 ~^ in11[2];
assign w1374 = in11[2] & w1248;
assign w1375 = in11[2] ~| w1248;
assign w1376 = w1249;
assign w1377 = w1130 ~^ w1250;
assign w1378 = w1130 | w1250;
assign w1379 = w1130 & w1250;
assign w1380 = w1131 ~^ w1251;
assign w1381 = w1129 ~^ w1252;
assign w1382 = w1129 | w1252;
assign w1383 = w1129 & w1252;
assign w1384 = w1124 | w1253;
assign w1385 = w578 ~^ w1254;
assign w1386 = w914 | w1254;
assign w1387 = w891 & w1255;
assign w1388 = w1244 ~^ w1256;
assign w1389 = w1119 | w1258;
assign w1390 = w902 ~^ w1261;
assign w1391 = w1096 | w1263;
assign w1392 = w925 ~^ w1264;
assign w1393 = w916 & w1265;
assign w1394 = w904 ~^ w1267;
assign w1395 = w904 ~| w1268;
assign w1396 = w620 ~^ w1269;
assign w1397 = w622 ~| w1269;
assign w1398 = w907 ~^ w1271;
assign w1399 = w907 ~| w1272;
assign w1400 = w903 ~| w1274;
assign w1401 = w901 ~^ w1276;
assign w1402 = w901 ~| w1277;
assign w1403 = w1137 & w1279;
assign w1404 = ~w1280;
assign w1405 = w976 ~^ w1282;
assign w1406 = w1146 | w1282;
assign w1407 = w974 ~^ w1284;
assign w1408 = w1144 | w1284;
assign w1409 = w978 ~^ w1286;
assign w1410 = ~w1288;
assign w1411 = ~w1297;
assign w1412 = w1168 & w1298;
assign w1413 = w1171 & w1300;
assign w1414 = w1174 & w1302;
assign w1415 = ~w1303;
assign w1416 = w1178 & w1304;
assign w1417 = ~w1305;
assign w1418 = ~w1306;
assign w1419 = w1182 & w1307;
assign w1420 = w1186 & w1309;
assign w1421 = ~w1310;
assign w1422 = ~w1312;
assign w1423 = w1196 & w1315;
assign w1424 = w1199 & w1316;
assign w1425 = w1201 & w1317;
assign w1426 = w1229 ~| w1318;
assign w1427 = w1066 ~^ w1319;
assign w1428 = w1067 | w1319;
assign w1429 = w1209 & w1320;
assign w1430 = w1218 & w1322;
assign w1431 = w1222 & w1323;
assign w1432 = w1034 ~^ w1324;
assign w1433 = w1034 | w1325;
assign w1434 = w1040 | w1326;
assign w1435 = w1014 ~^ w1327;
assign w1436 = w989 | w1328;
assign w1437 = w989 & w1328;
assign w1438 = w1020 ~^ w1329;
assign w1439 = w1020 | w1330;
assign w1440 = w986 | w1331;
assign w1441 = w1044 ~^ w1332;
assign w1442 = w1044 | w1333;
assign w1443 = in3[28] | w1334;
assign w1444 = w1004 ~^ w1335;
assign w1445 = w1004 | w1336;
assign w1446 = in3[24] | w1337;
assign w1447 = w1203 | w1339;
assign w1448 = w1018 ~^ w1340;
assign w1449 = w1018 | w1341;
assign w1450 = w987 | w1342;
assign w1451 = w1156 ~^ w1343;
assign w1452 = w1287 ~| w1343;
assign w1453 = ~w1343;
assign w1454 = w1050 | w1344;
assign w1455 = w1030 | w1345;
assign w1456 = ~w1346;
assign w1457 = w1005 ~^ w1347;
assign w1458 = w686 | w1348;
assign w1459 = w1005 | w1349;
assign w1460 = ~w1350;
assign w1461 = w181 | w1351;
assign w1462 = w1013 ~^ w1352;
assign w1463 = w1013 | w1353;
assign w1464 = w994 | w1354;
assign w1465 = w1022 ~^ w1355;
assign w1466 = w1022 | w1356;
assign w1467 = in3[26] | w1357;
assign w1468 = w1016 ~^ w1358;
assign w1469 = w991 | w1359;
assign w1470 = w1016 | w1360;
assign w1471 = ~w1361;
assign w1472 = w1153 ~| w1362;
assign w1473 = ~w1362;
assign w1474 = w1138 ~^ w1363;
assign w1475 = w1138 | w1364;
assign w1476 = w1043 | w1365;
assign w1477 = w1368;
assign w1478 = w1121 | w1369;
assign w1479 = ~w1369;
assign w1480 = w912 ~^ w1370;
assign w1481 = w1106 | w1371;
assign w1482 = w1367 ~^ w1373;
assign w1483 = w1367 ~| w1375;
assign w1484 = w238 ~| w1376;
assign w1485 = w909 ~^ w1377;
assign w1486 = w1105 | w1379;
assign w1487 = w903 ~^ w1380;
assign w1488 = w908 ~^ w1381;
assign w1489 = w1104 | w1383;
assign w1490 = w1124 ~^ w1385;
assign w1491 = w1384 & w1386;
assign w1492 = w1387;
assign w1493 = w1388;
assign w1494 = w1244 & w1389;
assign w1495 = w1262 & w1391;
assign w1496 = w1122 ~^ w1393;
assign w1497 = w1259 ~| w1393;
assign w1498 = w939 ~^ w1394;
assign w1499 = ~w1394;
assign w1500 = w918 | w1395;
assign w1501 = w221 ~| w1396;
assign w1502 = w621 | w1397;
assign w1503 = w931 ~^ w1398;
assign w1504 = ~w1398;
assign w1505 = w920 | w1399;
assign w1506 = w1251 | w1400;
assign w1507 = w932 ~^ w1401;
assign w1508 = ~w1401;
assign w1509 = w919 | w1402;
assign w1510 = w1362 ~^ w1409;
assign w1511 = w1361 ~| w1411;
assign w1512 = w1306 ~^ w1412;
assign w1513 = ~w1413;
assign w1514 = w1297 ~^ w1414;
assign w1515 = w1312 ~^ w1416;
assign w1516 = w1346 ~| w1417;
assign w1517 = w1303 ~^ w1419;
assign w1518 = w1404 ~^ w1420;
assign w1519 = w1280 ~| w1420;
assign w1520 = ~w1420;
assign w1521 = w1219 ~^ w1423;
assign w1522 = w1221 | w1423;
assign w1523 = w1308 | w1424;
assign w1524 = w1308 & w1424;
assign w1525 = w1403 ~^ w1424;
assign w1526 = w1311 ~^ w1425;
assign w1527 = ~w1427;
assign w1528 = w1068 & w1428;
assign w1529 = w1010 ~^ w1429;
assign w1530 = w1010 | w1429;
assign w1531 = w1010 & w1429;
assign w1532 = w1305 ~^ w1430;
assign w1533 = w1310 ~^ w1431;
assign w1534 = w1295 ~| w1432;
assign w1535 = ~w1432;
assign w1536 = w1433 & w1434;
assign w1537 = w1422 ~| w1435;
assign w1538 = ~w1435;
assign w1539 = w1014 | w1437;
assign w1540 = w1418 ~| w1438;
assign w1541 = ~w1438;
assign w1542 = w1439 & w1440;
assign w1543 = w1442 & w1443;
assign w1544 = w1410 ~^ w1444;
assign w1545 = w1410 ~| w1444;
assign w1546 = ~w1444;
assign w1547 = w1445 & w1446;
assign w1548 = ~w1448;
assign w1549 = w1449 & w1450;
assign w1550 = w1156 | w1453;
assign w1551 = w1454 & w1455;
assign w1552 = w1305 | w1456;
assign w1553 = w1421 ~| w1457;
assign w1554 = ~w1457;
assign w1555 = w1458 & w1459;
assign w1556 = w1441 ~^ w1461;
assign w1557 = w1441 ~| w1461;
assign w1558 = w1441 & w1461;
assign w1559 = w1415 ~| w1462;
assign w1560 = ~w1462;
assign w1561 = w1463 & w1464;
assign w1562 = ~w1465;
assign w1563 = w1466 & w1467;
assign w1564 = w1469 & w1470;
assign w1565 = w1297 | w1471;
assign w1566 = w1150 | w1472;
assign w1567 = w1286 | w1473;
assign w1568 = ~w1474;
assign w1569 = w1475 & w1476;
assign w1570 = w239 ~| w1477;
assign w1571 = w1390 & w1478;
assign w1572 = w937 ~^ w1479;
assign w1573 = w937 ~| w1479;
assign w1574 = w938 ~^ w1480;
assign w1575 = ~w1480;
assign w1576 = w1372 & w1481;
assign w1577 = ~w1482;
assign w1578 = w1374 | w1483;
assign w1579 = w866 ~| w1484;
assign w1580 = w940 ~^ w1485;
assign w1581 = ~w1485;
assign w1582 = w1378 & w1486;
assign w1583 = w936 ~^ w1487;
assign w1584 = ~w1487;
assign w1585 = w941 ~^ w1488;
assign w1586 = ~w1488;
assign w1587 = w1382 & w1489;
assign w1588 = w945 ~^ w1490;
assign w1589 = ~w1490;
assign w1590 = w1392 ~^ w1491;
assign w1591 = w1112 & w1491;
assign w1592 = w1112 ~| w1491;
assign w1593 = w1492 ~^ in11[3];
assign w1594 = in11[3] | w1492;
assign w1595 = in11[3] & w1492;
assign w1596 = w884 & w1493;
assign w1597 = w1257 | w1494;
assign w1598 = w1496;
assign w1599 = w1260 | w1497;
assign w1600 = w939 ~| w1499;
assign w1601 = w939 & w1499;
assign w1602 = w1266 & w1500;
assign w1603 = w853 ~| w1501;
assign w1604 = w1502;
assign w1605 = w931 ~| w1504;
assign w1606 = w931 & w1504;
assign w1607 = w1270 & w1505;
assign w1608 = w1273 & w1506;
assign w1609 = w932 & w1508;
assign w1610 = w932 ~| w1508;
assign w1611 = w1275 & w1509;
assign w1612 = ~w1510;
assign w1613 = w1414 | w1511;
assign w1614 = w1438 ~^ w1512;
assign w1615 = w1361 ~^ w1514;
assign w1616 = w1435 ~^ w1515;
assign w1617 = w1430 | w1516;
assign w1618 = w1462 ~^ w1517;
assign w1619 = w1468 ~^ w1518;
assign w1620 = w1404 | w1520;
assign w1621 = w1301 | w1521;
assign w1622 = w1301 & w1521;
assign w1623 = w1220 & w1522;
assign w1624 = w1403 | w1524;
assign w1625 = w1308 ~^ w1525;
assign w1626 = w1448 ~^ w1526;
assign w1627 = w187 ~^ w1528;
assign w1628 = w341 & w1528;
assign w1629 = w341 ~| w1528;
assign w1630 = w1346 ~^ w1532;
assign w1631 = w1457 ^ w1533;
assign w1632 = w1164 | w1535;
assign w1633 = w1053 ~^ w1536;
assign w1634 = w1053 & w1536;
assign w1635 = w1053 ~| w1536;
assign w1636 = w1416 | w1537;
assign w1637 = w1312 | w1538;
assign w1638 = w1436 & w1539;
assign w1639 = w1412 | w1540;
assign w1640 = w1306 | w1541;
assign w1641 = w1407 ~^ w1542;
assign w1642 = w1283 | w1542;
assign w1643 = w1338 ~^ w1543;
assign w1644 = w1426 | w1543;
assign w1645 = w1288 | w1546;
assign w1646 = w1534 | w1547;
assign w1647 = w1295 ^ w1547;
assign w1648 = w1311 | w1548;
assign w1649 = w1311 & w1548;
assign w1650 = w1289 ~^ w1549;
assign w1651 = w1290 | w1549;
assign w1652 = w1213 ~^ w1551;
assign w1653 = w1215 | w1551;
assign w1654 = w1431 | w1553;
assign w1655 = w1310 | w1554;
assign w1656 = w1292 ~^ w1555;
assign w1657 = w1294 | w1555;
assign w1658 = w1419 | w1559;
assign w1659 = w1303 | w1560;
assign w1660 = w1405 ~^ w1561;
assign w1661 = w1281 | w1561;
assign w1662 = w1206 ~^ w1563;
assign w1663 = w1207 | w1563;
assign w1664 = w1529 ~^ w1564;
assign w1665 = w1531 | w1564;
assign w1666 = w1566 & w1567;
assign w1667 = w1313 ~^ w1569;
assign w1668 = w1313 | w1569;
assign w1669 = w1313 & w1569;
assign w1670 = w875 ~| w1570;
assign w1671 = w1390 ~^ w1572;
assign w1672 = w1571 | w1573;
assign w1673 = w938 ~| w1575;
assign w1674 = w938 & w1575;
assign w1675 = w940 & w1581;
assign w1676 = w940 ~| w1581;
assign w1677 = w1574 ~^ w1582;
assign w1678 = w936 ~| w1584;
assign w1679 = w936 & w1584;
assign w1680 = w1495 ~^ w1585;
assign w1681 = w941 ~| w1586;
assign w1682 = w941 & w1586;
assign w1683 = w1583 ~^ w1587;
assign w1684 = w1576 ~^ w1588;
assign w1685 = w945 & w1589;
assign w1686 = w945 ~| w1589;
assign w1687 = w1590;
assign w1688 = w1264 ~| w1591;
assign w1689 = w1596;
assign w1690 = w1597;
assign w1691 = w898 & w1598;
assign w1692 = w1599;
assign w1693 = w1507 ~^ w1602;
assign w1694 = w892 & w1604;
assign w1695 = w1498 ~^ w1607;
assign w1696 = w1601 ~| w1607;
assign w1697 = w1503 ~^ w1608;
assign w1698 = w1606 ~| w1608;
assign w1699 = w1602 ~| w1609;
assign w1700 = w1580 ~^ w1611;
assign w1701 = w1565 & w1613;
assign w1702 = ~w1614;
assign w1703 = ~w1615;
assign w1704 = w1552 & w1617;
assign w1705 = ~w1618;
assign w1706 = ~w1619;
assign w1707 = w1468 & w1620;
assign w1708 = ~w1623;
assign w1709 = w1523 & w1624;
assign w1710 = ~w1625;
assign w1711 = ~w1626;
assign w1712 = ~w1630;
assign w1713 = w1296 ~^ w1633;
assign w1714 = w1296 ~| w1634;
assign w1715 = w1636 & w1637;
assign w1716 = w1147 ~^ w1638;
assign w1717 = w1149 | w1638;
assign w1718 = w1639 & w1640;
assign w1719 = ~w1641;
assign w1720 = w1408 & w1642;
assign w1721 = ~w1643;
assign w1722 = w1447 & w1644;
assign w1723 = w1632 & w1646;
assign w1724 = w1432 ~^ w1647;
assign w1725 = w1425 | w1649;
assign w1726 = w1291 & w1651;
assign w1727 = ~w1652;
assign w1728 = w1214 & w1653;
assign w1729 = w1654 & w1655;
assign w1730 = w1293 & w1657;
assign w1731 = w1658 & w1659;
assign w1732 = ~w1660;
assign w1733 = w1406 & w1661;
assign w1734 = w1350 ~^ w1662;
assign w1735 = w1460 ~| w1662;
assign w1736 = ~w1662;
assign w1737 = w1208 & w1663;
assign w1738 = w1451 ~^ w1664;
assign w1739 = w1452 | w1664;
assign w1740 = w1530 & w1665;
assign w1741 = ~w1666;
assign w1742 = w1671;
assign w1743 = w1672;
assign w1744 = w1582 ~| w1674;
assign w1745 = w1611 ~| w1675;
assign w1746 = w1677;
assign w1747 = w1587 ~| w1679;
assign w1748 = w1680;
assign w1749 = w1495 ~| w1682;
assign w1750 = w1683;
assign w1751 = w1684;
assign w1752 = w1576 ~| w1685;
assign w1753 = w900 & w1687;
assign w1754 = w1592 | w1688;
assign w1755 = w1689 ~^ in11[4];
assign w1756 = w220 ~| w1690;
assign w1757 = w1691 ~^ in11[15];
assign w1758 = w895 & w1692;
assign w1759 = w1693;
assign w1760 = ~w1694;
assign w1761 = w1695;
assign w1762 = w1600 | w1696;
assign w1763 = w1697;
assign w1764 = w1605 | w1698;
assign w1765 = w1610 | w1699;
assign w1766 = w1700;
assign w1767 = w1519 | w1707;
assign w1768 = w1667 ~^ w1709;
assign w1769 = w1669 | w1709;
assign w1770 = w1562 | w1713;
assign w1771 = ~w1713;
assign w1772 = w1635 | w1714;
assign w1773 = w1148 & w1717;
assign w1774 = w1666 | w1719;
assign w1775 = w1660 ~^ w1720;
assign w1776 = ~w1720;
assign w1777 = w1527 ~^ w1722;
assign w1778 = w1427 | w1722;
assign w1779 = ~w1722;
assign w1780 = ~w1724;
assign w1781 = w1648 & w1725;
assign w1782 = w1656 ~^ w1726;
assign w1783 = w1656 | w1726;
assign w1784 = w1656 & w1726;
assign w1785 = w1724 ~^ w1728;
assign w1786 = ~w1728;
assign w1787 = w1474 ~^ w1730;
assign w1788 = w1568 | w1730;
assign w1789 = ~w1730;
assign w1790 = w1720 | w1732;
assign w1791 = w1716 ~^ w1733;
assign w1792 = w1716 | w1733;
assign w1793 = w1716 & w1733;
assign w1794 = w1350 | w1736;
assign w1795 = w1556 ~^ w1737;
assign w1796 = w1557 ~| w1737;
assign w1797 = ~w1738;
assign w1798 = w1550 & w1739;
assign w1799 = w1544 ~^ w1740;
assign w1800 = w1545 | w1740;
assign w1801 = w1641 ~^ w1741;
assign w1802 = w1641 ~| w1741;
assign w1803 = w896 & w1742;
assign w1804 = w242 ~| w1743;
assign w1805 = w1673 | w1744;
assign w1806 = w1676 | w1745;
assign w1807 = w893 & w1746;
assign w1808 = w1678 | w1747;
assign w1809 = w889 & w1748;
assign w1810 = w1681 | w1749;
assign w1811 = w888 & w1750;
assign w1812 = w894 & w1751;
assign w1813 = w1686 | w1752;
assign w1814 = w1753;
assign w1815 = w1754;
assign w1816 = w871 ~| w1756;
assign w1817 = ~w1758;
assign w1818 = w887 & w1759;
assign w1819 = w886 & w1761;
assign w1820 = w1762;
assign w1821 = w885 & w1763;
assign w1822 = w1764;
assign w1823 = w1765;
assign w1824 = w897 & w1766;
assign w1825 = w1738 ~| w1767;
assign w1826 = ~w1767;
assign w1827 = w1619 | w1768;
assign w1828 = ~w1768;
assign w1829 = w1668 & w1769;
assign w1830 = w1465 ~^ w1771;
assign w1831 = w1465 ~| w1771;
assign w1832 = w1734 ~^ w1772;
assign w1833 = w1650 | w1773;
assign w1834 = w1650 & w1773;
assign w1835 = w1731 ~^ w1775;
assign w1836 = w1660 ~| w1776;
assign w1837 = w1527 ~| w1779;
assign w1838 = w1728 | w1780;
assign w1839 = w1773 ~^ w1781;
assign w1840 = w1729 ~^ w1782;
assign w1841 = w1729 | w1784;
assign w1842 = w1724 ~| w1786;
assign w1843 = w1704 ~^ w1787;
assign w1844 = w1474 ~| w1789;
assign w1845 = w1715 ~^ w1791;
assign w1846 = w1715 | w1793;
assign w1847 = w1772 & w1794;
assign w1848 = ~w1795;
assign w1849 = w1558 | w1796;
assign w1850 = w1652 | w1799;
assign w1851 = ~w1799;
assign w1852 = w1645 & w1800;
assign w1853 = w1718 ~^ w1801;
assign w1854 = w1718 | w1802;
assign w1855 = w1803 ~^ in11[5];
assign w1856 = w870 ~| w1804;
assign w1857 = w1805;
assign w1858 = w1806;
assign w1859 = w1807 ~^ in11[12];
assign w1860 = w1808;
assign w1861 = w1809;
assign w1862 = w1810;
assign w1863 = w1811;
assign w1864 = w1812 ~^ in11[13];
assign w1865 = w1813;
assign w1866 = w1814 ~^ in11[14];
assign w1867 = in11[14] & w1814;
assign w1868 = in11[14] | w1814;
assign w1869 = w242 ~| w1815;
assign w1870 = w1818;
assign w1871 = w1819;
assign w1872 = w216 ~| w1820;
assign w1873 = w1821;
assign w1874 = w244 ~| w1822;
assign w1875 = w241 ~| w1823;
assign w1876 = w1824;
assign w1877 = w1738 ~^ w1826;
assign w1878 = w1797 | w1826;
assign w1879 = w1706 ~^ w1828;
assign w1880 = w1706 ~| w1828;
assign w1881 = w1825 | w1829;
assign w1882 = w1723 ~^ w1830;
assign w1883 = w1723 | w1831;
assign w1884 = ~w1832;
assign w1885 = w1781 | w1834;
assign w1886 = w1616 ~^ w1835;
assign w1887 = w1616 & w1835;
assign w1888 = w1616 ~| w1835;
assign w1889 = w1731 | w1836;
assign w1890 = w1650 ~^ w1839;
assign w1891 = w1712 | w1840;
assign w1892 = ~w1840;
assign w1893 = w1783 & w1841;
assign w1894 = w1710 ~^ w1843;
assign w1895 = w1710 ~| w1843;
assign w1896 = ~w1843;
assign w1897 = w1704 | w1844;
assign w1898 = w1626 ~^ w1845;
assign w1899 = w1711 | w1845;
assign w1900 = ~w1845;
assign w1901 = w1792 & w1846;
assign w1902 = w1735 | w1847;
assign w1903 = w1643 ~| w1849;
assign w1904 = ~w1849;
assign w1905 = w1652 ~^ w1851;
assign w1906 = w1727 ~| w1851;
assign w1907 = w1785 ~^ w1852;
assign w1908 = w1842 | w1852;
assign w1909 = w1618 ^ w1853;
assign w1910 = w1774 & w1854;
assign w1911 = w220 ~| w1857;
assign w1912 = w240 ~| w1858;
assign w1913 = w240 ~| w1860;
assign w1914 = w1861 ~^ in11[6];
assign w1915 = w216 ~| w1862;
assign w1916 = w1863 ~^ in11[7];
assign w1917 = w215 ~| w1865;
assign w1918 = w854 ~| w1869;
assign w1919 = w1870 ~^ in11[10];
assign w1920 = in11[10] & w1870;
assign w1921 = in11[10] | w1870;
assign w1922 = w1871 ~^ in11[9];
assign w1923 = in11[9] & w1871;
assign w1924 = in11[9] | w1871;
assign w1925 = w851 ~| w1872;
assign w1926 = w1873 ~^ in11[8];
assign w1927 = in11[8] | w1873;
assign w1928 = in11[8] & w1873;
assign w1929 = w877 ~| w1874;
assign w1930 = w856 ~| w1875;
assign w1931 = w1876 ~^ in11[11];
assign w1932 = in11[11] & w1876;
assign w1933 = in11[11] | w1876;
assign w1934 = w1829 ^ w1877;
assign w1935 = w1878 & w1881;
assign w1936 = ~w1882;
assign w1937 = w1770 & w1883;
assign w1938 = w1833 & w1885;
assign w1939 = w1790 & w1889;
assign w1940 = w1631 | w1890;
assign w1941 = w1631 & w1890;
assign w1942 = w1630 ~| w1892;
assign w1943 = w1893 ~^ w1894;
assign w1944 = w1893 | w1895;
assign w1945 = w1625 | w1896;
assign w1946 = w1788 & w1897;
assign w1947 = w1626 ~| w1900;
assign w1948 = w1631 ^ w1901;
assign w1949 = w1795 ~^ w1902;
assign w1950 = w1848 ~| w1902;
assign w1951 = ~w1902;
assign w1952 = w1643 ~^ w1904;
assign w1953 = w1721 | w1904;
assign w1954 = w1798 ~^ w1905;
assign w1955 = w1798 | w1906;
assign w1956 = ~w1907;
assign w1957 = w1838 & w1908;
assign w1958 = w1886 ~^ w1910;
assign w1959 = w1888 ~| w1910;
assign w1960 = w864 ~| w1911;
assign w1961 = w874 ~| w1912;
assign w1962 = w869 ~| w1913;
assign w1963 = w880 ~| w1915;
assign w1964 = w876 ~| w1917;
assign w1965 = ~w1934;
assign w1966 = w1884 ~^ w1937;
assign w1967 = w1832 | w1937;
assign w1968 = ~w1937;
assign w1969 = w1630 ~^ w1938;
assign w1970 = w1898 ~^ w1939;
assign w1971 = w1901 | w1941;
assign w1972 = w1938 | w1942;
assign w1973 = ~w1943;
assign w1974 = w1944 & w1945;
assign w1975 = w1879 ~^ w1946;
assign w1976 = w1880 | w1946;
assign w1977 = w1939 | w1947;
assign w1978 = w1890 ~^ w1948;
assign w1979 = w1795 | w1951;
assign w1980 = w1935 ~^ w1954;
assign w1981 = ~w1954;
assign w1982 = w1850 & w1955;
assign w1983 = w1936 ~^ w1957;
assign w1984 = w1882 | w1957;
assign w1985 = ~w1957;
assign w1986 = ~w1958;
assign w1987 = w1887 | w1959;
assign w1988 = w1884 ~| w1968;
assign w1989 = w1840 ~^ w1969;
assign w1990 = ~w1970;
assign w1991 = w1940 & w1971;
assign w1992 = w1891 & w1972;
assign w1993 = ~w1974;
assign w1994 = w1974 | w1975;
assign w1995 = ~w1975;
assign w1996 = w1827 & w1976;
assign w1997 = w1899 & w1977;
assign w1998 = ~w1978;
assign w1999 = w1935 | w1981;
assign w2000 = w1935 & w1981;
assign w2001 = w1907 ~^ w1982;
assign w2002 = w1956 | w1982;
assign w2003 = w1956 & w1982;
assign w2004 = w1936 ~| w1985;
assign w2005 = w1970 ~| w1987;
assign w2006 = ~w1987;
assign w2007 = ~w1989;
assign w2008 = w1989 ~^ w1991;
assign w2009 = ~w1991;
assign w2010 = w1973 ~^ w1992;
assign w2011 = w1943 | w1992;
assign w2012 = ~w1992;
assign w2013 = w1974 ~^ w1995;
assign w2014 = w1993 ~| w1995;
assign w2015 = w1965 ~^ w1996;
assign w2016 = w1934 | w1996;
assign w2017 = ~w1996;
assign w2018 = w1978 ~^ w1997;
assign w2019 = ~w1997;
assign w2020 = w1997 | w1998;
assign w2021 = w1970 ~^ w2006;
assign w2022 = w1990 | w2006;
assign w2023 = w1991 | w2007;
assign w2024 = w1989 ~| w2009;
assign w2025 = w1973 ~| w2012;
assign w2026 = w1965 ~| w2017;
assign w2027 = w1978 ~| w2019;
wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027;
endmodule
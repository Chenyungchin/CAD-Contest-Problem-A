module top(in1, in2, in3, in4, out1);
input wire [15:0] in1;
input wire [15:0] in2;
input wire [15:0] in3;
input wire [1:0] in4;
output wire [31:0] out1;
assign or = ~in4[0];
assign or = in1[5] & in4[1];
assign or = in1[3] & in4[1];
assign or = in1[2] & in4[1];
assign or = in1[4] & in4[1];
assign or = in1[7] & in4[1];
assign or = in1[0] & in4[1];
assign or = in1[8] & in4[1];
assign or = in1[15] & in4[1];
assign or = in1[1] & in4[1];
assign or = in1[14] & in4[1];
assign or = in1[13] & in4[1];
assign or = in1[12] & in4[1];
assign or = in1[6] & in4[1];
assign or = in1[10] & in4[1];
assign or = in1[9] & in4[1];
assign or = in1[11] & in4[1];
assign and = in4[1] | in4[0];
assign and = ~in4[1];
assign and = ~in4[1];
assign and = ~in4[1];
assign and = ~in4[1];
assign and = ~in4[1];
assign and = ~in4[1];
assign and = ~in4[1];
assign and = ~in4[1];
assign and = ~in4[1];
endmodule
module top(in1, in2, in3, in4, out1);
input wire [15:0] in1;
input wire [15:0] in2;
input wire [15:0] in3;
input wire [15:0] in4;
output wire [33:0] out1;
assign w0 = ~in1[0];
assign w1 = ~in1[1];
assign w2 = in1[2] ~| in1[0];
assign w3 = ~in1[2];
assign w4 = in1[3] ~^ in1[1];
assign w5 = ~in1[3];
assign w6 = ~in1[4];
assign w7 = ~in1[5];
assign w8 = ~in1[6];
assign w9 = in1[7] ~^ in1[2];
assign w10 = ~in1[7];
assign w11 = in1[8] ~^ in1[6];
assign w12 = in1[8] | in1[6];
assign w13 = ~in1[8];
assign w14 = in1[9] ~^ in1[4];
assign w15 = ~in1[9];
assign w16 = in1[10] ~^ in1[5];
assign w17 = ~in1[10];
assign w18 = in1[11] ~^ in1[6];
assign w19 = ~in1[11];
assign w20 = in1[12] ~^ in1[7];
assign w21 = ~in1[12];
assign w22 = in1[13] ~^ in1[8];
assign w23 = ~in1[13];
assign w24 = ~in1[14];
assign w25 = ~in1[15];
assign w26 = in1[6] ~| in2[0];
assign w27 = in1[6] & in2[0];
assign w28 = ~in2[0];
assign w29 = in1[2] ~^ in2[1];
assign w30 = ~in2[1];
assign w31 = ~in2[2];
assign w32 = ~in2[4];
assign w33 = ~in2[5];
assign w34 = in2[6] ~^ in2[3];
assign w35 = ~in2[6];
assign w36 = in2[8] ~^ in2[5];
assign w37 = in2[9] ~^ in2[6];
assign w38 = ~in2[9];
assign w39 = in2[10] ~^ in2[7];
assign w40 = in1[14] ~| in2[10];
assign w41 = ~in2[10];
assign w42 = in2[11] ~^ in2[8];
assign w43 = in1[13] ~^ in2[11];
assign w44 = ~in2[11];
assign w45 = in2[12] ~^ in2[9];
assign w46 = ~in2[12];
assign w47 = in1[15] ~^ in2[13];
assign w48 = in1[15] ~| in2[13];
assign w49 = ~in2[13];
assign w50 = in1[10] ~^ in2[14];
assign w51 = in1[10] ~| in2[14];
assign w52 = ~in2[14];
assign w53 = in2[15] ~^ in2[12];
assign w54 = ~in2[15];
assign w55 = ~in3[0];
assign w56 = ~in3[2];
assign w57 = ~in3[3];
assign w58 = ~in3[4];
assign w59 = ~in3[6];
assign w60 = ~in3[7];
assign w61 = ~in3[8];
assign w62 = ~in3[10];
assign w63 = ~in3[15];
assign w64 = in4[0] ~^ in3[0];
assign w65 = in4[0] ~^ in2[2];
assign w66 = in4[0] ~^ in1[4];
assign w67 = in4[0] ~^ in2[0];
assign w68 = ~in4[0];
assign w69 = in4[1] ~^ in3[1];
assign w70 = ~in4[1];
assign w71 = in4[2] ~^ in2[2];
assign w72 = in4[2] ~^ in2[7];
assign w73 = in4[2] ~^ in3[2];
assign w74 = in4[2] ~| in2[7];
assign w75 = in4[2] ~| in4[0];
assign w76 = in4[2] & in2[7];
assign w77 = ~in4[2];
assign w78 = in4[3] ~^ in1[5];
assign w79 = in4[3] ~^ in2[3];
assign w80 = in4[3] ~^ in2[4];
assign w81 = in4[3] ~^ in3[3];
assign w82 = in4[3] ~| in2[4];
assign w83 = ~in4[3];
assign w84 = in4[4] ~^ in1[4];
assign w85 = in4[4] ~^ in2[4];
assign w86 = in4[4] ~^ in1[1];
assign w87 = in4[4] ~^ in3[4];
assign w88 = in4[4] ~| in1[1];
assign w89 = ~in4[4];
assign w90 = in4[5] ~^ in1[7];
assign w91 = in4[5] ~^ in3[5];
assign w92 = in4[5] ~^ in2[5];
assign w93 = in4[5] | in4[1];
assign w94 = ~in4[5];
assign w95 = in4[6] ~^ in1[8];
assign w96 = in4[6] ~^ in2[6];
assign w97 = in4[6] ~^ in3[6];
assign w98 = in4[6] ~| in4[0];
assign w99 = in4[6] ~| in4[2];
assign w100 = ~in4[6];
assign w101 = in4[7] ~| in2[6];
assign w102 = ~in4[7];
assign w103 = in4[8] ~^ in4[1];
assign w104 = in4[8] ~^ in3[8];
assign w105 = in4[8] & in1[9];
assign w106 = in4[8] ~| in4[1];
assign w107 = in4[8] | in1[9];
assign w108 = ~in4[8];
assign w109 = in4[9] ~^ in3[9];
assign w110 = in4[9] ~| in2[8];
assign w111 = in4[9] | in4[5];
assign w112 = in4[9] & in2[8];
assign w113 = in4[9] ~| in2[15];
assign w114 = ~in4[9];
assign w115 = in4[10] ~^ in2[13];
assign w116 = in4[10] ~^ in3[10];
assign w117 = in4[10] ~| in2[9];
assign w118 = ~in4[10];
assign w119 = in4[11] ~^ in3[11];
assign w120 = in4[11] ~| in2[10];
assign w121 = in4[11] | in4[7];
assign w122 = in4[11] & in4[7];
assign w123 = in4[11] & in2[10];
assign w124 = ~in4[11];
assign w125 = in4[12] ~^ in4[11];
assign w126 = in4[12] ~^ in3[12];
assign w127 = in4[12] | in4[8];
assign w128 = in4[12] ~| in2[11];
assign w129 = in4[12] & in4[8];
assign w130 = in4[12] ~| in4[11];
assign w131 = in4[12] & in2[11];
assign w132 = ~in4[12];
assign w133 = in4[13] ~^ in4[12];
assign w134 = in4[13] ~^ in3[13];
assign w135 = in4[13] ~| in2[12];
assign w136 = in4[13] & in4[9];
assign w137 = in4[13] | in4[9];
assign w138 = ~in4[13];
assign w139 = in4[14] ~^ in4[12];
assign w140 = in4[14] ~^ in4[10];
assign w141 = in4[14] ~^ in3[14];
assign w142 = in4[14] ~^ in4[13];
assign w143 = in4[14] & in4[12];
assign w144 = in4[14] ~| in4[12];
assign w145 = in4[14] | in4[10];
assign w146 = in4[14] & in4[10];
assign w147 = ~in4[14];
assign w148 = in4[15] ~^ in4[11];
assign w149 = in4[15] ~^ in3[15];
assign w150 = in4[15] ~^ in4[13];
assign w151 = in4[15] ~^ in4[14];
assign w152 = in4[15] ~^ in2[15];
assign w153 = ~in4[15];
assign  = 1'b0;
assign w154 = w0 ~| in4[0];
assign w155 = w1 | in4[1];
assign w156 = in4[1] & w1;
assign w157 = w0 | w3;
assign w158 = w4 ~^ in4[1];
assign w159 = w6 | in4[4];
assign w160 = in4[4] & w6;
assign w161 = w7 ~| in4[3];
assign w162 = w9 ~^ in4[1];
assign w163 = w10 ~| in4[5];
assign w164 = w10 | in4[1];
assign w165 = w13 ~| in4[6];
assign w166 = w8 ~| w13;
assign w167 = w14 ~^ in4[3];
assign w168 = w15 | in4[0];
assign w169 = w15 ~| in4[3];
assign w170 = w16 ~^ in4[4];
assign w171 = w17 ~| in4[4];
assign w172 = w18 ~^ in4[5];
assign w173 = w19 | in4[2];
assign w174 = w19 ~| in4[5];
assign w175 = in4[2] & w19;
assign w176 = w20 ~^ in4[6];
assign w177 = in4[3] & w21;
assign w178 = w21 | in4[3];
assign w179 = w21 | in4[6];
assign w180 = w22 ~^ in4[7];
assign w181 = w23 | in4[7];
assign w182 = w23 | in4[4];
assign w183 = w24 | in2[15];
assign w184 = w24 | in4[5];
assign w185 = w25 ~| in4[6];
assign w186 = w25 | in4[9];
assign w187 = w26 | w27;
assign w188 = ~w27;
assign w189 = ~w27;
assign w190 = in1[2] & w30;
assign w191 = w30 | in1[2];
assign w192 = w34 ~^ in4[7];
assign w193 = w36 ~^ in4[9];
assign w194 = w37 ~^ in4[10];
assign w195 = w39 ~^ in4[11];
assign w196 = w39 ~^ in1[14];
assign w197 = w24 | w41;
assign w198 = w42 ~^ in4[8];
assign w199 = w42 ~^ in4[12];
assign w200 = ~w43;
assign w201 = w44 | in4[8];
assign w202 = w23 & w44;
assign w203 = w45 ~^ in4[13];
assign w204 = w49 | in4[10];
assign w205 = w25 ~| w49;
assign w206 = w17 | w52;
assign w207 = w53 ~^ in4[9];
assign w208 = w53 ~^ in1[14];
assign w209 = w54 ~| in1[14];
assign out1[0] = w64 ~^ in1[0];
assign w210 = w65 ~^ in4[6];
assign w211 = w66 ~^ in4[2];
assign w212 = w67 ~^ in1[9];
assign w213 = w68 | in1[0];
assign w214 = w68 ~| in1[9];
assign w215 = w69 ~^ in1[1];
assign w216 = w70 ~| in1[7];
assign w217 = w71 ~^ in1[11];
assign w218 = w72 ~^ in2[4];
assign w219 = w73 ~^ in4[0];
assign w220 = w68 ~| w73;
assign w221 = ~w73;
assign w222 = in2[4] ~| w74;
assign w223 = in1[4] | w75;
assign w224 = w68 | w77;
assign w225 = w56 | w77;
assign w226 = w78 ~^ in1[3];
assign w227 = w79 ~^ in1[12];
assign w228 = w80 ~^ in2[1];
assign w229 = w81 ~^ in2[0];
assign w230 = in2[1] | w82;
assign w231 = w83 | in1[5];
assign w232 = w57 | w83;
assign w233 = w83 | in1[9];
assign w234 = w32 | w83;
assign w235 = w84 ~^ in2[3];
assign w236 = w85 ~^ in1[13];
assign w237 = w86 ~^ in2[5];
assign w238 = w33 ~| w88;
assign w239 = w89 ~| in1[13];
assign w240 = w89 | in1[10];
assign w241 = w58 | w89;
assign w242 = w1 ~| w89;
assign w243 = w90 ~^ in1[5];
assign w244 = w91 ~^ in4[1];
assign w245 = w92 ~^ in1[14];
assign w246 = in3[5] & w93;
assign w247 = w94 ~| in1[14];
assign w248 = w70 ~| w94;
assign w249 = w94 | in1[7];
assign w250 = w94 | in1[11];
assign w251 = w95 ~^ in1[3];
assign w252 = w96 ~^ in1[15];
assign w253 = w97 ~^ in4[2];
assign w254 = in2[2] | w98;
assign w255 = w59 | w99;
assign w256 = w100 | in1[15];
assign w257 = w100 ~| in1[12];
assign w258 = w100 | in1[8];
assign w259 = w68 | w100;
assign w260 = w77 | w100;
assign w261 = in2[3] | w101;
assign w262 = w102 ~^ in3[7];
assign w263 = w102 ~| in1[13];
assign w264 = w35 | w102;
assign w265 = w60 | w102;
assign w266 = w103 ~^ in2[1];
assign w267 = w11 ~^ w104;
assign w268 = w30 ~| w106;
assign w269 = ~w107;
assign w270 = w108 ~| in2[11];
assign w271 = w70 ~| w108;
assign w272 = w61 | w108;
assign w273 = w109 ~^ in4[5];
assign w274 = in2[5] ~| w110;
assign w275 = in3[9] & w111;
assign w276 = in2[12] | w113;
assign w277 = w114 | in1[15];
assign w278 = w54 | w114;
assign w279 = w94 ~| w114;
assign w280 = w115 ~^ in2[10];
assign w281 = w116 ~^ in1[10];
assign w282 = in1[10] ~| w116;
assign w283 = ~w116;
assign w284 = in2[6] ~| w117;
assign w285 = w118 ~| in2[13];
assign w286 = w38 ~| w118;
assign w287 = w62 | w118;
assign w288 = w119 ~^ in4[7];
assign w289 = in2[7] ~| w120;
assign w290 = in3[11] & w121;
assign w291 = w125 ~^ in2[14];
assign w292 = w126 ~^ in4[8];
assign w293 = in3[12] & w127;
assign w294 = in2[8] ~| w128;
assign w295 = in2[14] | w130;
assign w296 = w124 | w132;
assign w297 = ~w133;
assign w298 = w134 ~^ in4[9];
assign w299 = in2[9] | w135;
assign w300 = in3[13] & w137;
assign w301 = w46 | w138;
assign w302 = w132 | w138;
assign w303 = w139 ~^ in4[7];
assign w304 = w140 ~^ in1[11];
assign w305 = w141 ~^ in4[10];
assign w306 = w102 ~| w144;
assign w307 = in3[14] & w145;
assign w308 = ~w145;
assign w309 = w138 | w147;
assign w310 = w148 ~^ in1[12];
assign w311 = w149 ~^ in4[11];
assign w312 = w50 ~^ w150;
assign w313 = w51 | w150;
assign w314 = ~w152;
assign w315 = w124 & w153;
assign w316 = w147 & w153;
assign w317 = w124 | w153;
assign w318 = w138 | w153;
assign w319 = w54 & w153;
assign w320 = in3[0] | w154;
assign w321 = in3[1] & w155;
assign w322 = ~w155;
assign w323 = ~w156;
assign w324 = ~w157;
assign w325 = w157 ~^ w158;
assign w326 = w157 | w158;
assign w327 = in2[3] & w159;
assign w328 = in1[3] | w161;
assign w329 = ~w162;
assign w330 = in1[5] | w163;
assign w331 = in1[2] & w164;
assign w332 = w5 | w165;
assign w333 = w104 | w166;
assign w334 = in2[0] & w168;
assign w335 = w6 | w169;
assign w336 = w7 | w171;
assign w337 = in2[2] & w173;
assign w338 = w8 | w174;
assign w339 = in2[3] & w178;
assign w340 = in1[7] & w179;
assign w341 = ~w180;
assign w342 = in1[8] & w181;
assign w343 = in2[4] & w182;
assign w344 = in2[5] & w184;
assign w345 = w35 | w185;
assign w346 = ~w187;
assign w347 = ~w193;
assign w348 = w170 & w194;
assign w349 = w170 | w194;
assign w350 = w172 | w195;
assign w351 = w172 & w195;
assign w352 = in2[7] & w197;
assign w353 = w176 | w199;
assign w354 = w176 & w199;
assign w355 = in2[8] & w201;
assign w356 = w133 ~| w202;
assign w357 = ~w202;
assign w358 = w180 ~| w203;
assign w359 = ~w203;
assign w360 = in2[10] & w204;
assign w361 = w46 | w209;
assign w362 = ~w210;
assign w363 = w87 | w211;
assign w364 = w87 & w211;
assign w365 = w215 ~^ in3[0];
assign w366 = w55 | w215;
assign w367 = w55 & w215;
assign w368 = w167 | w217;
assign w369 = w167 & w217;
assign w370 = in4[0] | w221;
assign w371 = w76 | w222;
assign w372 = w223 & w224;
assign w373 = w28 & w225;
assign w374 = w28 | w225;
assign w375 = ~w227;
assign w376 = ~w228;
assign w377 = w225 ~^ w229;
assign w378 = w29 ~^ w232;
assign w379 = w190 | w232;
assign w380 = w230 & w234;
assign w381 = ~w235;
assign w382 = ~w236;
assign w383 = w210 ~^ w237;
assign w384 = ~w237;
assign w385 = w241 ~^ in2[2];
assign w386 = w31 | w241;
assign w387 = w31 & w241;
assign w388 = w238 | w242;
assign w389 = w188 ~| w243;
assign w390 = w189 & w243;
assign w391 = w226 ~^ w244;
assign w392 = w226 & w244;
assign w393 = w226 ~| w244;
assign w394 = ~w245;
assign w395 = w246 | w248;
assign w396 = ~w251;
assign w397 = ~w252;
assign w398 = w235 ~^ w253;
assign w399 = ~w253;
assign w400 = w254 & w259;
assign w401 = w255 & w260;
assign w402 = in1[0] | w262;
assign w403 = ~w262;
assign w404 = w261 & w264;
assign w405 = w218 ~^ w266;
assign w406 = ~w266;
assign w407 = w105 | w269;
assign w408 = w268 | w271;
assign w409 = ~w272;
assign w410 = w162 ~^ w273;
assign w411 = ~w273;
assign w412 = w112 | w274;
assign w413 = w186 & w277;
assign w414 = w276 & w278;
assign w415 = w275 | w279;
assign w416 = ~w280;
assign w417 = w17 | w283;
assign w418 = w284 | w286;
assign w419 = ~w287;
assign w420 = w193 ~^ w288;
assign w421 = ~w288;
assign w422 = w123 | w289;
assign w423 = w122 | w290;
assign w424 = ~w291;
assign w425 = w227 ~^ w292;
assign w426 = ~w292;
assign w427 = w129 | w293;
assign w428 = w131 | w294;
assign w429 = w295 & w296;
assign w430 = w236 ~^ w298;
assign w431 = ~w298;
assign w432 = w136 | w300;
assign w433 = w299 & w301;
assign w434 = w47 ~^ w302;
assign w435 = w48 ~| w302;
assign w436 = w196 ~^ w303;
assign w437 = w196 & w303;
assign w438 = w196 | w303;
assign w439 = w186 ~^ w304;
assign w440 = w186 & w304;
assign w441 = w186 ~| w304;
assign w442 = w245 ~^ w305;
assign w443 = ~w305;
assign w444 = w143 | w306;
assign w445 = w146 | w307;
assign w446 = w19 ~| w308;
assign w447 = w309 ~^ in2[14];
assign w448 = w52 ~| w309;
assign w449 = ~w309;
assign w450 = w280 ~^ w310;
assign w451 = ~w310;
assign w452 = w252 ~^ w311;
assign w453 = w206 & w313;
assign w454 = w63 | w315;
assign w455 = w21 ~| w315;
assign w456 = w152 ~^ w316;
assign w457 = w314 ~| w316;
assign w458 = ~w316;
assign w459 = ~w317;
assign w460 = w318 ~^ in2[9];
assign w461 = w38 ~| w318;
assign w462 = ~w318;
assign w463 = w213 & w320;
assign w464 = w156 | w321;
assign w465 = in1[3] | w322;
assign w466 = w2 | w324;
assign w467 = ~w324;
assign w468 = w160 | w327;
assign w469 = w231 & w328;
assign w470 = w273 ~| w329;
assign w471 = w249 & w330;
assign w472 = w216 | w331;
assign w473 = w258 & w332;
assign w474 = w12 & w333;
assign w475 = w214 | w334;
assign w476 = w233 & w335;
assign w477 = w240 & w336;
assign w478 = w175 | w337;
assign w479 = w250 & w338;
assign w480 = w177 | w339;
assign w481 = w257 | w340;
assign w482 = w263 | w342;
assign w483 = w239 | w343;
assign w484 = w247 | w344;
assign w485 = w256 & w345;
assign w486 = w288 ~| w347;
assign w487 = w40 | w352;
assign w488 = w270 | w355;
assign w489 = w297 | w357;
assign w490 = w341 | w359;
assign w491 = w285 | w360;
assign w492 = w183 & w361;
assign w493 = w237 ~| w362;
assign w494 = w81 | w373;
assign w495 = w292 | w375;
assign w496 = ~w378;
assign w497 = w191 & w379;
assign w498 = w253 ~| w381;
assign w499 = w298 | w382;
assign w500 = w267 ~^ w383;
assign w501 = w210 | w384;
assign w502 = w372 ^ w385;
assign w503 = w372 | w387;
assign w504 = ~w388;
assign w505 = w305 | w394;
assign w506 = w266 ~| w396;
assign w507 = w311 | w397;
assign w508 = w311 & w397;
assign w509 = w235 | w399;
assign w510 = w272 | w400;
assign w511 = ~w400;
assign w512 = w389 ~| w401;
assign w513 = w189 ^ w401;
assign w514 = w403 ~^ in1[0];
assign w515 = w0 ~| w403;
assign w516 = w251 ~^ w405;
assign w517 = w251 | w406;
assign w518 = ~w407;
assign w519 = w287 ~^ w408;
assign w520 = ~w408;
assign w521 = w212 ~^ w410;
assign w522 = w162 | w411;
assign w523 = w198 ~^ w413;
assign w524 = w312 | w413;
assign w525 = w312 & w413;
assign w526 = ~w414;
assign w527 = ~w415;
assign w528 = w310 | w416;
assign w529 = ~w418;
assign w530 = w408 | w419;
assign w531 = w193 | w421;
assign w532 = w227 ~| w426;
assign w533 = ~w428;
assign w534 = w208 ~^ w429;
assign w535 = w236 ~| w431;
assign w536 = w142 & w434;
assign w537 = w142 | w434;
assign w538 = w205 | w435;
assign w539 = w207 ~^ w439;
assign w540 = w207 ~| w441;
assign w541 = w245 ~| w443;
assign w542 = w146 | w446;
assign w543 = w151 ~^ w447;
assign w544 = in2[14] | w449;
assign w545 = w280 ~| w451;
assign w546 = ~w453;
assign w547 = w317 & w454;
assign w548 = w152 | w458;
assign w549 = w455 | w459;
assign w550 = in2[9] | w462;
assign out1[1] = w365 ~^ w463;
assign w551 = w367 | w463;
assign w552 = w219 ~^ w464;
assign w553 = w370 & w464;
assign w554 = w323 & w465;
assign w555 = ~w466;
assign w556 = w158 & w467;
assign w557 = w402 & w468;
assign w558 = w395 ~^ w469;
assign w559 = w346 ~| w469;
assign w560 = ~w469;
assign w561 = w212 | w470;
assign w562 = w265 ~^ w471;
assign w563 = w265 | w471;
assign w564 = w265 & w471;
assign w565 = w415 ~^ w472;
assign w566 = w415 ~| w472;
assign w567 = ~w472;
assign w568 = w369 | w473;
assign w569 = w217 ^ w473;
assign w570 = w192 ~^ w474;
assign w571 = w192 | w474;
assign w572 = w192 & w474;
assign w573 = w281 ~^ w475;
assign w574 = w417 & w475;
assign w575 = w348 | w476;
assign w576 = w170 ^ w476;
assign w577 = w351 | w477;
assign w578 = w172 ^ w477;
assign w579 = w412 ~^ w478;
assign w580 = w412 | w478;
assign w581 = w412 & w478;
assign w582 = w354 | w479;
assign w583 = w176 ^ w479;
assign w584 = w418 | w480;
assign w585 = ~w480;
assign w586 = w180 ~^ w481;
assign w587 = in2[13] ~| w482;
assign w588 = in2[13] & w482;
assign w589 = w422 ~^ w483;
assign w590 = w422 & w483;
assign w591 = w422 | w483;
assign w592 = w428 | w484;
assign w593 = ~w484;
assign w594 = w433 ~^ w485;
assign w595 = w107 | w487;
assign w596 = ~w487;
assign w597 = w460 ~^ w488;
assign w598 = ~w489;
assign w599 = w481 & w490;
assign w600 = w424 | w491;
assign w601 = w424 & w491;
assign w602 = w142 ^ w492;
assign w603 = w267 | w493;
assign w604 = w374 & w494;
assign w605 = w391 ~^ w497;
assign w606 = w393 ~| w497;
assign w607 = ~w500;
assign w608 = w386 & w503;
assign w609 = w218 | w506;
assign w610 = w272 ~^ w511;
assign w611 = w409 ~| w511;
assign w612 = w390 | w512;
assign w613 = w243 ~^ w513;
assign w614 = w468 ~^ w514;
assign w615 = ~w516;
assign w616 = w485 ~| w518;
assign w617 = w485 & w518;
assign w618 = w371 ~^ w519;
assign w619 = w287 ~| w520;
assign w620 = ~w521;
assign w621 = w312 ~^ w523;
assign w622 = w198 | w525;
assign w623 = w480 ~^ w529;
assign w624 = w371 & w530;
assign w625 = w484 ~^ w533;
assign w626 = w492 | w536;
assign w627 = ~w538;
assign w628 = w440 | w540;
assign w629 = w526 & w542;
assign w630 = ~w542;
assign w631 = w538 ~^ w543;
assign w632 = ~w543;
assign w633 = w151 & w544;
assign w634 = w547 ^ in2[13];
assign w635 = w491 ~^ w549;
assign w636 = w488 & w550;
assign w637 = w366 & w551;
assign w638 = w466 ~^ w552;
assign w639 = w220 | w553;
assign w640 = w364 | w554;
assign w641 = w87 ~^ w554;
assign w642 = w552 & w555;
assign w643 = w552 ~| w555;
assign w644 = w515 | w557;
assign w645 = w187 ~^ w558;
assign w646 = w187 | w560;
assign w647 = w522 & w561;
assign w648 = w380 ^ w562;
assign w649 = w380 | w564;
assign w650 = w404 ~^ w565;
assign w651 = w404 | w566;
assign w652 = w527 | w567;
assign w653 = w368 & w568;
assign w654 = w167 ~^ w569;
assign w655 = ~w573;
assign w656 = w282 | w574;
assign w657 = w349 & w575;
assign w658 = w194 ~^ w576;
assign w659 = w350 & w577;
assign w660 = w195 ~^ w578;
assign w661 = w423 ~^ w579;
assign w662 = w423 & w580;
assign w663 = w353 & w582;
assign w664 = w199 ~^ w583;
assign w665 = w427 & w584;
assign w666 = w529 ~| w585;
assign w667 = w203 ~^ w586;
assign w668 = w547 ~| w587;
assign w669 = w432 ~^ w589;
assign w670 = w432 & w591;
assign w671 = w445 & w592;
assign w672 = w533 ~| w593;
assign w673 = w407 ~^ w594;
assign w674 = w444 & w595;
assign w675 = w444 ~^ w596;
assign w676 = w269 ~| w596;
assign w677 = w453 ~| w597;
assign w678 = ~w597;
assign w679 = w356 | w598;
assign w680 = ~w598;
assign w681 = w358 | w599;
assign w682 = w549 & w600;
assign w683 = w434 ~^ w602;
assign w684 = w501 & w603;
assign w685 = w378 ~^ w604;
assign w686 = w496 | w604;
assign w687 = w496 & w604;
assign w688 = w502 & w605;
assign w689 = w502 | w605;
assign w690 = w392 | w606;
assign w691 = w398 ~^ w608;
assign w692 = w498 | w608;
assign w693 = w517 & w609;
assign w694 = w388 ~^ w610;
assign w695 = w504 | w611;
assign w696 = ~w613;
assign w697 = w228 ~^ w614;
assign w698 = w228 ~| w614;
assign w699 = ~w614;
assign w700 = w433 ~| w617;
assign w701 = ~w621;
assign w702 = w524 & w622;
assign w703 = w427 ~^ w623;
assign w704 = w619 | w624;
assign w705 = w445 ~^ w625;
assign w706 = w537 & w626;
assign w707 = w543 | w627;
assign w708 = w414 & w630;
assign w709 = w538 ~| w632;
assign w710 = w448 | w633;
assign w711 = w482 ~^ w634;
assign w712 = w291 ~^ w635;
assign w713 = w461 | w636;
assign out1[2] = w637 ~^ w638;
assign w714 = w325 ~^ w639;
assign w715 = w326 & w639;
assign w716 = w363 & w640;
assign w717 = w211 ~^ w641;
assign w718 = w637 ~| w642;
assign w719 = ~w645;
assign w720 = w395 & w646;
assign w721 = w516 ~^ w647;
assign w722 = w644 ~^ w648;
assign w723 = w644 & w648;
assign w724 = w644 | w648;
assign w725 = w563 & w649;
assign w726 = ~w650;
assign w727 = w651 & w652;
assign w728 = ~w654;
assign w729 = w650 | w655;
assign w730 = ~w656;
assign w731 = ~w658;
assign w732 = ~w660;
assign w733 = w658 ~| w661;
assign w734 = ~w661;
assign w735 = w581 | w662;
assign w736 = ~w664;
assign w737 = w665 | w666;
assign w738 = ~w667;
assign w739 = w588 | w668;
assign w740 = w664 ~| w669;
assign w741 = ~w669;
assign w742 = w590 | w670;
assign w743 = w671 | w672;
assign w744 = w107 ^ w675;
assign w745 = w674 | w676;
assign w746 = w546 | w678;
assign w747 = w534 ~^ w679;
assign w748 = ~w679;
assign w749 = w673 ~^ w681;
assign w750 = ~w681;
assign w751 = w601 | w682;
assign w752 = w489 ~^ w683;
assign w753 = w680 & w683;
assign w754 = w489 | w683;
assign w755 = w645 ~^ w690;
assign w756 = ~w690;
assign w757 = ~w691;
assign w758 = w509 & w692;
assign w759 = w656 ~^ w693;
assign w760 = w620 | w694;
assign w761 = ~w694;
assign w762 = w510 & w695;
assign w763 = w376 | w699;
assign w764 = w616 | w700;
assign w765 = w539 ~^ w702;
assign w766 = w539 | w702;
assign w767 = w539 & w702;
assign w768 = ~w703;
assign w769 = w425 ~^ w704;
assign w770 = w495 & w704;
assign w771 = ~w705;
assign w772 = w631 ~^ w706;
assign w773 = w43 ~^ w708;
assign w774 = w629 | w708;
assign w775 = ~w708;
assign w776 = w706 | w709;
assign w777 = w456 ~^ w710;
assign w778 = w548 & w710;
assign w779 = w673 & w711;
assign w780 = w673 ~| w711;
assign w781 = w450 ~^ w713;
assign w782 = w528 & w713;
assign w783 = w377 ~^ w714;
assign w784 = w377 & w714;
assign w785 = w377 | w714;
assign w786 = w556 | w715;
assign w787 = w688 | w716;
assign w788 = w502 ^ w716;
assign w789 = w685 ~^ w717;
assign w790 = w687 | w717;
assign w791 = w643 | w718;
assign w792 = w690 ~| w719;
assign w793 = w559 | w720;
assign w794 = w612 ~^ w722;
assign w795 = w612 & w724;
assign w796 = w570 ~^ w725;
assign w797 = w572 | w725;
assign w798 = w573 ~| w726;
assign w799 = w486 | w727;
assign w800 = w420 ^ w727;
assign w801 = w618 | w730;
assign w802 = w618 & w730;
assign w803 = w703 | w732;
assign w804 = w653 | w733;
assign w805 = w731 | w734;
assign w806 = w653 ~^ w734;
assign w807 = w430 ~^ w735;
assign w808 = w499 & w735;
assign w809 = w442 ~^ w737;
assign w810 = w505 & w737;
assign w811 = w705 | w738;
assign w812 = w659 | w740;
assign w813 = w736 | w741;
assign w814 = w659 ~^ w741;
assign w815 = w452 ~^ w742;
assign w816 = w507 & w742;
assign w817 = w436 ~^ w743;
assign w818 = w438 & w743;
assign w819 = ~w744;
assign w820 = w453 ~^ w745;
assign w821 = w745 & w746;
assign w822 = ~w747;
assign w823 = w208 & w748;
assign w824 = w208 ~| w748;
assign w825 = w711 ~^ w749;
assign w826 = w747 ~| w751;
assign w827 = ~w751;
assign w828 = w691 ~^ w755;
assign w829 = w645 | w756;
assign w830 = w613 ~^ w758;
assign w831 = w696 ~| w758;
assign w832 = ~w758;
assign w833 = w618 ~^ w759;
assign w834 = w521 ~^ w761;
assign w835 = w521 ~| w761;
assign w836 = w655 ^ w762;
assign w837 = w744 | w764;
assign w838 = ~w764;
assign w839 = w660 ~| w768;
assign w840 = w657 ~^ w768;
assign w841 = ~w769;
assign w842 = w532 | w770;
assign w843 = w667 ~| w771;
assign w844 = w663 ~^ w771;
assign w845 = w712 ~^ w773;
assign w846 = w628 ~^ w774;
assign w847 = w628 | w774;
assign w848 = w628 & w774;
assign w849 = w43 ~| w775;
assign w850 = ~w775;
assign w851 = w707 & w776;
assign w852 = ~w777;
assign w853 = w457 | w778;
assign w854 = w750 ~| w780;
assign w855 = w545 | w782;
assign w856 = ~w786;
assign w857 = w689 & w787;
assign w858 = w605 ~^ w788;
assign w859 = w786 ~^ w789;
assign w860 = w786 ~| w789;
assign w861 = ~w789;
assign w862 = w686 & w790;
assign out1[3] = w783 ~^ w791;
assign w863 = w785 & w791;
assign w864 = w757 | w792;
assign w865 = w697 ~^ w793;
assign w866 = w763 & w793;
assign w867 = ~w794;
assign w868 = w723 | w795;
assign w869 = ~w796;
assign w870 = w571 & w797;
assign w871 = w762 | w798;
assign w872 = w531 & w799;
assign w873 = w654 ~^ w800;
assign w874 = w728 ~| w800;
assign w875 = w728 & w800;
assign w876 = w693 | w802;
assign w877 = w804 & w805;
assign w878 = w658 ~^ w806;
assign w879 = ~w807;
assign w880 = w535 | w808;
assign w881 = ~w809;
assign w882 = w541 | w810;
assign w883 = w812 & w813;
assign w884 = w664 ~^ w814;
assign w885 = ~w815;
assign w886 = w508 | w816;
assign w887 = ~w817;
assign w888 = w437 | w818;
assign w889 = w597 ~^ w820;
assign w890 = w677 | w821;
assign w891 = w751 ~^ w822;
assign w892 = w429 ~| w823;
assign w893 = ~w825;
assign w894 = w822 | w827;
assign w895 = w613 | w832;
assign w896 = ~w833;
assign w897 = w684 ~^ w834;
assign w898 = w684 | w835;
assign w899 = w726 ~^ w836;
assign w900 = w739 & w837;
assign w901 = w819 ~| w838;
assign w902 = w739 ~^ w838;
assign w903 = w657 | w839;
assign w904 = w660 ~^ w840;
assign w905 = w807 ~^ w842;
assign w906 = ~w842;
assign w907 = w663 | w843;
assign w908 = w667 ~^ w844;
assign w909 = w712 | w849;
assign w910 = w200 | w850;
assign w911 = w777 ~^ w851;
assign w912 = ~w851;
assign w913 = ~w852;
assign w914 = w319 ~^ w853;
assign w915 = w319 | w853;
assign w916 = w319 & w853;
assign w917 = w779 | w854;
assign w918 = w845 ~^ w855;
assign w919 = w845 & w855;
assign w920 = w845 | w855;
assign w921 = w828 ~^ w857;
assign w922 = w828 | w857;
assign w923 = w828 & w857;
assign w924 = ~w858;
assign w925 = w856 | w861;
assign w926 = w858 ~^ w862;
assign w927 = w784 | w863;
assign w928 = w829 & w864;
assign w929 = w830 ~^ w865;
assign w930 = w698 | w866;
assign w931 = ~w868;
assign w932 = w868 ~^ w869;
assign w933 = w868 ~| w869;
assign w934 = w615 | w870;
assign w935 = ~w870;
assign w936 = w729 & w871;
assign w937 = w769 | w872;
assign w938 = ~w872;
assign w939 = w801 & w876;
assign w940 = ~w878;
assign w941 = w842 ~| w879;
assign w942 = w809 ~^ w880;
assign w943 = ~w880;
assign w944 = w880 ~| w881;
assign w945 = w815 ~^ w882;
assign w946 = ~w882;
assign w947 = ~w884;
assign w948 = w882 ~| w885;
assign w949 = w817 ~^ w886;
assign w950 = w817 ~| w886;
assign w951 = ~w886;
assign w952 = w621 ~^ w888;
assign w953 = w701 ~| w888;
assign w954 = ~w888;
assign w955 = ~w889;
assign w956 = w846 ~^ w890;
assign w957 = w847 & w890;
assign w958 = w824 | w892;
assign w959 = w865 & w895;
assign w960 = w760 & w898;
assign w961 = ~w899;
assign w962 = w900 | w901;
assign w963 = w819 ~^ w902;
assign w964 = w803 & w903;
assign w965 = ~w904;
assign w966 = w877 ^ w905;
assign w967 = w807 | w906;
assign w968 = w811 & w907;
assign w969 = w909 & w910;
assign w970 = w852 | w912;
assign w971 = w851 ~| w913;
assign w972 = ~w917;
assign w973 = w862 ~| w924;
assign w974 = w862 & w924;
assign out1[4] = w859 ~^ w927;
assign w975 = ~w927;
assign w976 = ~w928;
assign w977 = w928 | w929;
assign w978 = ~w929;
assign w979 = w500 ~| w930;
assign w980 = ~w930;
assign w981 = w796 | w931;
assign w982 = w897 ~^ w932;
assign w983 = w897 | w933;
assign w984 = w721 ~^ w935;
assign w985 = w516 ~| w935;
assign w986 = w873 ~^ w936;
assign w987 = w875 ~| w936;
assign w988 = w841 ~^ w938;
assign w989 = w841 ~| w938;
assign w990 = w877 | w941;
assign w991 = w809 | w943;
assign w992 = w883 ~^ w945;
assign w993 = w815 | w946;
assign w994 = w883 | w948;
assign w995 = w887 | w951;
assign w996 = w917 ~^ w952;
assign w997 = w621 | w954;
assign w998 = w781 ~^ w956;
assign w999 = ~w956;
assign w1000 = w848 | w957;
assign w1001 = w752 ~^ w958;
assign w1002 = w754 & w958;
assign w1003 = w831 | w959;
assign w1004 = w960 ~^ w961;
assign w1005 = w765 ~^ w962;
assign w1006 = ~w962;
assign w1007 = ~w963;
assign w1008 = w944 | w964;
assign w1009 = w942 ^ w964;
assign w1010 = w904 | w966;
assign w1011 = ~w966;
assign w1012 = w949 ~^ w968;
assign w1013 = w950 | w968;
assign w1014 = w891 ~^ w969;
assign w1015 = w826 | w969;
assign w1016 = w953 | w972;
assign w1017 = w860 | w975;
assign w1018 = w976 ~^ w978;
assign w1019 = w976 ~| w978;
assign w1020 = w867 | w979;
assign w1021 = w500 ~^ w980;
assign w1022 = w607 | w980;
assign w1023 = ~w982;
assign w1024 = w981 & w983;
assign w1025 = w899 | w984;
assign w1026 = ~w984;
assign w1027 = w647 | w985;
assign w1028 = ~w986;
assign w1029 = w874 | w987;
assign w1030 = w939 ~^ w988;
assign w1031 = w939 | w989;
assign w1032 = w967 & w990;
assign w1033 = w908 ~^ w992;
assign w1034 = ~w992;
assign w1035 = w993 & w994;
assign w1036 = ~w996;
assign w1037 = w781 & w999;
assign w1038 = w781 ~| w999;
assign w1039 = w918 ~^ w1000;
assign w1040 = w920 & w1000;
assign w1041 = ~w1001;
assign w1042 = w753 | w1002;
assign w1043 = ~w1003;
assign w1044 = w955 ~^ w1005;
assign w1045 = w889 ~| w1005;
assign w1046 = ~w1005;
assign w1047 = w767 | w1006;
assign w1048 = w996 | w1007;
assign w1049 = w991 & w1008;
assign w1050 = w947 | w1009;
assign w1051 = ~w1009;
assign w1052 = w965 ~| w1011;
assign w1053 = w893 | w1012;
assign w1054 = ~w1012;
assign w1055 = w995 & w1013;
assign w1056 = w894 & w1015;
assign w1057 = w997 & w1016;
assign w1058 = w925 & w1017;
assign w1059 = w794 ~^ w1021;
assign w1060 = w1020 & w1022;
assign w1061 = ~w1024;
assign w1062 = w1004 ~^ w1026;
assign w1063 = w961 ~| w1026;
assign w1064 = w934 & w1027;
assign w1065 = ~w1029;
assign w1066 = w940 | w1030;
assign w1067 = ~w1030;
assign w1068 = w937 & w1031;
assign w1069 = w908 | w1034;
assign w1070 = w908 & w1034;
assign w1071 = w1007 ~^ w1036;
assign w1072 = w963 ~| w1036;
assign w1073 = w919 | w1040;
assign w1074 = w772 ~^ w1042;
assign w1075 = w772 & w1042;
assign w1076 = w772 | w1042;
assign w1077 = w955 | w1046;
assign w1078 = w766 & w1047;
assign w1079 = w1033 ^ w1049;
assign w1080 = w947 ~^ w1051;
assign w1081 = w884 ~| w1051;
assign w1082 = w893 ~^ w1054;
assign w1083 = w825 ~| w1054;
assign w1084 = w1041 ~^ w1056;
assign w1085 = w1041 ~| w1056;
assign w1086 = ~w1056;
assign w1087 = w1045 | w1057;
assign w1088 = w1044 ^ w1057;
assign out1[5] = w926 ~^ w1058;
assign w1089 = w974 ~| w1058;
assign w1090 = w1043 | w1059;
assign w1091 = ~w1059;
assign w1092 = w982 | w1060;
assign w1093 = ~w1060;
assign w1094 = w1024 | w1062;
assign w1095 = ~w1062;
assign w1096 = w960 | w1063;
assign w1097 = w896 | w1064;
assign w1098 = ~w1064;
assign w1099 = w940 ~^ w1067;
assign w1100 = w878 ~| w1067;
assign w1101 = w1052 | w1068;
assign w1102 = w965 ~^ w1068;
assign w1103 = w1049 | w1070;
assign w1104 = w1055 ^ w1071;
assign w1105 = w1055 | w1072;
assign w1106 = w1014 ~^ w1073;
assign w1107 = w1014 | w1073;
assign w1108 = w1014 & w1073;
assign w1109 = w998 ~^ w1078;
assign w1110 = w1037 ~| w1078;
assign w1111 = ~w1079;
assign w1112 = w1032 ^ w1080;
assign w1113 = w1032 | w1081;
assign w1114 = w1035 ~^ w1082;
assign w1115 = w1035 | w1083;
assign w1116 = w1001 | w1086;
assign w1117 = w1077 & w1087;
assign w1118 = ~w1088;
assign w1119 = w973 | w1089;
assign w1120 = w1003 ~^ w1091;
assign w1121 = w1003 ~| w1091;
assign w1122 = w1023 ~^ w1093;
assign w1123 = w1023 ~| w1093;
assign w1124 = w1061 ~^ w1095;
assign w1125 = w1061 ~| w1095;
assign w1126 = w1025 & w1096;
assign w1127 = w896 ~^ w1098;
assign w1128 = w833 ~| w1098;
assign w1129 = w1029 ~^ w1099;
assign w1130 = w1065 | w1100;
assign w1131 = w1010 & w1101;
assign w1132 = w1011 ~^ w1102;
assign w1133 = w1069 & w1103;
assign w1134 = ~w1104;
assign w1135 = w1048 & w1105;
assign w1136 = ~w1109;
assign w1137 = w1038 | w1110;
assign w1138 = ~w1112;
assign w1139 = w1050 & w1113;
assign w1140 = ~w1114;
assign w1141 = w1053 & w1115;
assign w1142 = w1109 ~^ w1117;
assign out1[6] = w921 ~^ w1119;
assign w1143 = ~w1119;
assign w1144 = ~w1126;
assign w1145 = w986 ~^ w1127;
assign w1146 = w1028 | w1128;
assign w1147 = ~w1129;
assign w1148 = w1066 & w1130;
assign w1149 = w1112 | w1131;
assign w1150 = ~w1131;
assign w1151 = ~w1132;
assign w1152 = w1114 ~^ w1133;
assign w1153 = w1088 | w1135;
assign w1154 = ~w1135;
assign w1155 = w1117 ~| w1136;
assign w1156 = w1117 & w1136;
assign w1157 = w1039 ~^ w1137;
assign w1158 = w1039 & w1137;
assign w1159 = w1039 | w1137;
assign w1160 = w1131 ~^ w1138;
assign w1161 = w1079 | w1139;
assign w1162 = ~w1139;
assign w1163 = w1133 | w1140;
assign w1164 = w1133 & w1140;
assign w1165 = w1104 | w1141;
assign w1166 = ~w1141;
assign w1167 = w923 | w1143;
assign w1168 = w1126 | w1145;
assign w1169 = ~w1145;
assign w1170 = w1097 & w1146;
assign w1171 = w1132 | w1148;
assign w1172 = ~w1148;
assign w1173 = w1138 ~| w1150;
assign w1174 = w1118 ~^ w1154;
assign w1175 = w1118 ~| w1154;
assign w1176 = w1111 ~^ w1162;
assign w1177 = w1111 ~| w1162;
assign w1178 = w1134 ~^ w1166;
assign w1179 = w1134 ~| w1166;
assign w1180 = w922 & w1167;
assign w1181 = w1144 ~^ w1169;
assign w1182 = w1144 ~| w1169;
assign w1183 = w1129 | w1170;
assign w1184 = ~w1170;
assign w1185 = w1151 ~^ w1172;
assign w1186 = w1151 ~| w1172;
assign w1187 = w1019 | w1180;
assign out1[7] = w1018 ^ w1180;
assign w1188 = w1147 ~^ w1184;
assign w1189 = w1147 ~| w1184;
assign w1190 = w977 & w1187;
assign w1191 = w1121 | w1190;
assign out1[8] = w1120 ^ w1190;
assign w1192 = w1090 & w1191;
assign w1193 = w1123 | w1192;
assign out1[9] = w1122 ^ w1192;
assign w1194 = w1092 & w1193;
assign w1195 = w1125 | w1194;
assign out1[10] = w1124 ^ w1194;
assign w1196 = w1094 & w1195;
assign w1197 = w1182 | w1196;
assign out1[11] = w1181 ^ w1196;
assign w1198 = w1168 & w1197;
assign w1199 = w1189 | w1198;
assign out1[12] = w1188 ^ w1198;
assign w1200 = w1183 & w1199;
assign w1201 = w1186 | w1200;
assign out1[13] = w1185 ^ w1200;
assign w1202 = w1171 & w1201;
assign out1[14] = w1160 ~^ w1202;
assign w1203 = w1173 | w1202;
assign w1204 = w1149 & w1203;
assign w1205 = w1177 | w1204;
assign out1[15] = w1176 ^ w1204;
assign w1206 = w1161 & w1205;
assign out1[16] = w1152 ~^ w1206;
assign w1207 = w1164 | w1206;
assign w1208 = w1163 & w1207;
assign w1209 = w1179 | w1208;
assign out1[17] = w1178 ^ w1208;
assign w1210 = w1165 & w1209;
assign w1211 = w1175 | w1210;
assign out1[18] = w1174 ^ w1210;
assign w1212 = w1153 & w1211;
assign out1[19] = w1142 ~^ w1212;
assign w1213 = w1156 ~| w1212;
assign w1214 = w1155 | w1213;
assign out1[20] = w1157 ~^ w1214;
assign w1215 = w1159 & w1214;
assign w1216 = w1158 | w1215;
assign out1[21] = w1106 ~^ w1216;
assign w1217 = w1107 & w1216;
assign w1218 = w1108 | w1217;
assign out1[22] = w1084 ~^ w1218;
assign w1219 = w1116 & w1218;
assign w1220 = w1085 | w1219;
assign out1[23] = w1074 ~^ w1220;
assign w1221 = w1076 & w1220;
assign w1222 = w1075 | w1221;
assign out1[24] = w911 ~^ w1222;
assign w1223 = w970 & w1222;
assign w1224 = w971 | w1223;
assign out1[25] = w914 ~^ w1224;
assign w1225 = w915 & w1224;
assign w1226 = w916 ~| w1225;
assign out1[26] = w319 ~^ w1226;
wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226;
endmodule
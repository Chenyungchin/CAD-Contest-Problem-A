<<<<<<< HEAD
module top(a, b, ci, s, co);
input wire a;
input wire b;
input wire ci;
output wire co;
output wire s;
xnor g0(w0, a, b);
and g1(w1, a, b);
xnor g2(w2, w0, ci);
and g4(w3, ci, w0);
not g3(s, w2);
or g5(co, w1, w3);
wire w0, w1, w2, w3;
=======
module top(in1, in2, in3, out1);
input wire [3:0] in1;
input wire [3:0] in2;
input wire [3:0] in3;
output wire [3:0] out1;
assign w0 = ~in1[1];
assign w1 = in1[0] ~^ in2[0];
assign w2 = ~in2[1];
assign w3 = in1[2] | in2[2];
assign w4 = in1[2] & in2[2];
assign w5 = in3[0] & in2[0];
assign w6 = in3[0] | in2[0];
assign w7 = in3[1] ~^ in1[1];
assign w8 = ~in3[1];
assign w9 = in3[2] ~^ in2[2];
assign w10 = in3[3] ~^ in2[3];
assign out1[0] = w1 ~^ in3[0];
assign w11 = in3[2] & w3;
assign w12 = in1[0] & w6;
assign w13 = w7 ~^ in2[1];
assign w14 = w2 ~| w7;
assign w15 = ~w7;
assign w16 = w0 | w8;
assign w17 = w9 ~^ in1[2];
assign w18 = w10 ~^ in1[3];
assign w19 = w4 | w11;
assign w20 = w5 | w12;
assign w21 = in2[1] | w15;
assign w22 = ~w16;
assign w23 = w16 ~^ w17;
assign w24 = w18 ~^ w19;
assign out1[1] = w13 ^ w20;
assign w25 = w20 & w21;
assign w26 = w17 | w22;
assign w27 = w17 & w22;
assign w28 = w14 | w25;
assign out1[2] = w23 ^ w28;
assign w29 = w26 & w28;
assign w30 = w27 | w29;
assign out1[3] = w24 ~^ w30;
wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30;
>>>>>>> d1c140d2c15e97d61c0f2aece8dd425f3d8952b4
endmodule
module top(in1, in2, in3, in4, out1);
input wire [15:0] in1;
input wire [15:0] in2;
input wire [15:0] in3;
input wire [15:0] in4;
output wire [33:0] out1;
assign w0 = ~in1[0];
assign w1 = ~in1[1];
assign w2 = in1[2] ~| in1[0];
assign w3 = ~in1[2];
assign w4 = in1[3] ~^ in1[1];
assign w5 = ~in1[3];
assign w6 = ~in1[4];
assign w7 = ~in1[5];
assign w8 = ~in1[6];
assign w9 = in1[7] ~^ in1[2];
assign w10 = ~in1[7];
assign w11 = in1[8] ~^ in1[6];
assign w12 = in1[8] | in1[6];
assign w13 = ~in1[8];
assign w14 = in1[9] ~^ in1[4];
assign w15 = ~in1[9];
assign w16 = in1[10] ~^ in1[5];
assign w17 = ~in1[10];
assign w18 = in1[11] ~^ in1[6];
assign w19 = ~in1[11];
assign w20 = in1[12] ~^ in1[7];
assign w21 = ~in1[12];
assign w22 = in1[13] ~^ in1[8];
assign w23 = ~in1[13];
assign w24 = ~in1[14];
assign w25 = ~in1[15];
assign w26 = in1[6] ~| in2[0];
assign w27 = in1[6] & in2[0];
assign w28 = ~in2[0];
assign w29 = in1[2] ~^ in2[1];
assign w30 = ~in2[1];
assign w31 = ~in2[2];
assign w32 = ~in2[4];
assign w33 = ~in2[5];
assign w34 = in2[6] ~^ in2[3];
assign w35 = ~in2[6];
assign w36 = in2[8] ~^ in2[5];
assign w37 = in2[9] ~^ in2[6];
assign w38 = ~in2[9];
assign w39 = in2[10] ~^ in2[7];
assign w40 = in1[14] ~| in2[10];
assign w41 = ~in2[10];
assign w42 = in2[11] ~^ in2[8];
assign w43 = in1[13] ~^ in2[11];
assign w44 = ~in2[11];
assign w45 = in2[12] ~^ in2[9];
assign w46 = ~in2[12];
assign w47 = in1[15] ~^ in2[13];
assign w48 = in1[15] ~| in2[13];
assign w49 = ~in2[13];
assign w50 = in1[10] ~^ in2[14];
assign w51 = in1[10] ~| in2[14];
assign w52 = ~in2[14];
assign w53 = in2[15] ~^ in2[12];
assign w54 = ~in2[15];
assign w55 = ~in3[0];
assign w56 = ~in3[2];
assign w57 = ~in3[3];
assign w58 = ~in3[4];
assign w59 = ~in3[6];
assign w60 = ~in3[7];
assign w61 = ~in3[8];
assign w62 = ~in3[10];
assign w63 = ~in3[15];
assign w64 = in4[0] ~^ in3[0];
assign w65 = in4[0] ~^ in2[2];
assign w66 = in4[0] ~^ in1[4];
assign w67 = in4[0] ~^ in2[0];
assign w68 = ~in4[0];
assign w69 = in4[1] ~^ in3[1];
assign w70 = ~in4[1];
assign w71 = in4[2] ~^ in2[2];
assign w72 = in4[2] ~^ in2[7];
assign w73 = in4[2] ~^ in3[2];
assign w74 = in4[2] ~| in2[7];
assign w75 = in4[2] ~| in4[0];
assign w76 = in4[2] & in2[7];
assign w77 = ~in4[2];
assign w78 = in4[3] ~^ in1[5];
assign w79 = in4[3] ~^ in2[3];
assign w80 = in4[3] ~^ in2[4];
assign w81 = in4[3] ~^ in3[3];
assign w82 = in4[3] ~| in2[4];
assign w83 = ~in4[3];
assign w84 = in4[4] ~^ in1[4];
assign w85 = in4[4] ~^ in2[4];
assign w86 = in4[4] ~^ in1[1];
assign w87 = in4[4] ~^ in3[4];
assign w88 = in4[4] ~| in1[1];
assign w89 = ~in4[4];
assign w90 = in4[5] ~^ in1[7];
assign w91 = in4[5] ~^ in3[5];
assign w92 = in4[5] ~^ in2[5];
assign w93 = in4[5] | in4[1];
assign w94 = ~in4[5];
assign w95 = in4[6] ~^ in1[8];
assign w96 = in4[6] ~^ in2[6];
assign w97 = in4[6] ~^ in3[6];
assign w98 = in4[6] ~| in4[0];
assign w99 = in4[6] ~| in4[2];
assign w100 = ~in4[6];
assign w101 = in4[7] ~| in2[6];
assign w102 = ~in4[7];
assign w103 = in4[8] ~^ in4[1];
assign w104 = in4[8] ~^ in3[8];
assign w105 = in4[8] & in1[9];
assign w106 = in4[8] ~| in4[1];
assign w107 = in4[8] | in1[9];
assign w108 = ~in4[8];
assign w109 = in4[9] ~^ in3[9];
assign w110 = in4[9] ~| in2[8];
assign w111 = in4[9] | in4[5];
assign w112 = in4[9] & in2[8];
assign w113 = in4[9] ~| in2[15];
assign w114 = ~in4[9];
assign w115 = in4[10] ~^ in2[13];
assign w116 = in4[10] ~^ in3[10];
assign w117 = in4[10] ~| in2[9];
assign w118 = ~in4[10];
assign w119 = in4[11] ~^ in3[11];
assign w120 = in4[11] ~| in2[10];
assign w121 = in4[11] | in4[7];
assign w122 = in4[11] & in4[7];
assign w123 = in4[11] & in2[10];
assign w124 = ~in4[11];
assign w125 = in4[12] ~^ in4[11];
assign w126 = in4[12] ~^ in3[12];
assign w127 = in4[12] | in4[8];
assign w128 = in4[12] ~| in2[11];
assign w129 = in4[12] & in4[8];
assign w130 = in4[12] ~| in4[11];
assign w131 = in4[12] & in2[11];
assign w132 = ~in4[12];
assign w133 = in4[13] ~^ in4[12];
assign w134 = in4[13] ~^ in3[13];
assign w135 = in4[13] ~| in2[12];
assign w136 = in4[13] & in4[9];
assign w137 = in4[13] | in4[9];
assign w138 = ~in4[13];
assign w139 = in4[14] ~^ in4[12];
assign w140 = in4[14] ~^ in4[10];
assign w141 = in4[14] ~^ in3[14];
assign w142 = in4[14] ~^ in4[13];
assign w143 = in4[14] & in4[12];
assign w144 = in4[14] ~| in4[12];
assign w145 = in4[14] | in4[10];
assign w146 = in4[14] & in4[10];
assign w147 = ~in4[14];
assign w148 = in4[15] ~^ in4[11];
assign w149 = in4[15] ~^ in3[15];
assign w150 = in4[15] ~^ in4[13];
assign w151 = in4[15] ~^ in4[14];
assign w152 = in4[15] ~^ in2[15];
assign w153 = ~in4[15];

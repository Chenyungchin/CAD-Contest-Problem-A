module top(in1, in2, in3, out2);
input wire [31:0] in1;
input wire [31:0] in2;
input wire [31:0] in3;
output wire [40:0] out2;
assign w0 = ~in1[0];
assign w1 = ~in1[0];
assign w2 = ~in1[0];
assign w3 = ~in1[0];
assign w4 = ~in1[0];
assign w5 = ~in1[0];
assign w6 = ~in1[0];
assign w7 = ~in1[0];
assign w8 = ~in1[0];
assign w9 = ~in1[0];
assign w10 = ~in1[0];
assign w11 = ~in1[0];
assign w12 = ~in1[0];
assign w13 = ~in1[0];
assign w14 = ~in1[0];
assign w15 = ~in1[0];
assign w16 = in1[1] ~^ in1[0];
assign w17 = ~in1[1];
assign w18 = ~in1[1];
assign w19 = ~in1[1];
assign w20 = ~in1[1];
assign w21 = ~in1[1];
assign w22 = ~in1[1];
assign w23 = ~in1[1];
assign w24 = ~in1[1];
assign w25 = ~in1[1];
assign w26 = ~in1[1];
assign w27 = ~in1[1];
assign w28 = ~in1[1];
assign w29 = ~in1[1];
assign w30 = ~in1[1];
assign w31 = ~in1[1];
assign w32 = ~in1[1];
assign w33 = in1[2] ~^ in1[1];
assign w34 = ~in1[2];
assign w35 = ~in1[2];
assign w36 = ~in1[2];
assign w37 = ~in1[2];
assign w38 = ~in1[2];
assign w39 = ~in1[2];
assign w40 = ~in1[2];
assign w41 = ~in1[2];
assign w42 = ~in1[2];
assign w43 = ~in1[2];
assign w44 = ~in1[2];
assign w45 = ~in1[2];
assign w46 = ~in1[2];
assign w47 = ~in1[2];
assign w48 = ~in1[2];
assign w49 = ~in1[2];
assign w50 = in1[3] ~^ in1[2];
assign w51 = in1[3] ~| in1[2];
assign w52 = ~in1[3];
assign w53 = ~in1[3];
assign w54 = ~in1[3];
assign w55 = ~in1[3];
assign w56 = ~in1[3];
assign w57 = ~in1[3];
assign w58 = ~in1[3];
assign w59 = ~in1[3];
assign w60 = ~in1[3];
assign w61 = ~in1[3];
assign w62 = ~in1[3];
assign w63 = ~in1[3];
assign w64 = ~in1[3];
assign w65 = ~in1[3];
assign w66 = ~in1[3];
assign w67 = ~in1[3];
assign w68 = in1[4] ~^ in1[3];
assign w69 = in1[4] ~| in1[3];
assign w70 = ~in1[4];
assign w71 = ~in1[4];
assign w72 = ~in1[4];
assign w73 = ~in1[4];
assign w74 = ~in1[4];
assign w75 = ~in1[4];
assign w76 = ~in1[4];
assign w77 = ~in1[4];
assign w78 = ~in1[4];
assign w79 = ~in1[4];
assign w80 = ~in1[4];
assign w81 = ~in1[4];
assign w82 = ~in1[4];
assign w83 = ~in1[4];
assign w84 = ~in1[4];
assign w85 = ~in1[4];
assign w86 = in1[5] ~^ in1[4];
assign w87 = in1[5] ~| in1[4];
assign w88 = ~in1[5];
assign w89 = ~in1[5];
assign w90 = ~in1[5];
assign w91 = ~in1[5];
assign w92 = ~in1[5];
assign w93 = ~in1[5];
assign w94 = ~in1[5];
assign w95 = ~in1[5];
assign w96 = ~in1[5];
assign w97 = ~in1[5];
assign w98 = ~in1[5];
assign w99 = ~in1[5];
assign w100 = ~in1[5];
assign w101 = ~in1[5];
assign w102 = ~in1[5];
assign w103 = ~in1[5];
assign w104 = in1[6] ~^ in1[5];
assign w105 = in1[6] ~| in1[5];
assign w106 = ~in1[6];
assign w107 = ~in1[6];
assign w108 = ~in1[6];
assign w109 = ~in1[6];
assign w110 = ~in1[6];
assign w111 = ~in1[6];
assign w112 = ~in1[6];
assign w113 = ~in1[6];
assign w114 = ~in1[6];
assign w115 = ~in1[6];
assign w116 = ~in1[6];
assign w117 = ~in1[6];
assign w118 = ~in1[6];
assign w119 = ~in1[6];
assign w120 = ~in1[6];
assign w121 = ~in1[6];
assign w122 = in1[7] ~^ in1[6];
assign w123 = in1[7] ~| in1[6];
assign w124 = ~in1[7];
assign w125 = ~in1[7];
assign w126 = ~in1[7];
assign w127 = ~in1[7];
assign w128 = ~in1[7];
assign w129 = ~in1[7];
assign w130 = ~in1[7];
assign w131 = ~in1[7];
assign w132 = ~in1[7];
assign w133 = ~in1[7];
assign w134 = ~in1[7];
assign w135 = ~in1[7];
assign w136 = ~in1[7];
assign w137 = ~in1[7];
assign w138 = ~in1[7];
assign w139 = ~in1[7];
assign w140 = in1[8] ~^ in1[7];
assign w141 = in1[8] ~| in1[7];
assign w142 = ~in1[8];
assign w143 = ~in1[8];
assign w144 = ~in1[8];
assign w145 = ~in1[8];
assign w146 = ~in1[8];
assign w147 = ~in1[8];
assign w148 = ~in1[8];
assign w149 = ~in1[8];
assign w150 = ~in1[8];
assign w151 = ~in1[8];
assign w152 = ~in1[8];
assign w153 = ~in1[8];
assign w154 = ~in1[8];
assign w155 = ~in1[8];
assign w156 = ~in1[8];
assign w157 = ~in1[8];
assign w158 = in1[9] ~^ in1[8];
assign w159 = in1[9] ~| in1[8];
assign w160 = ~in1[9];
assign w161 = ~in1[9];
assign w162 = ~in1[9];
assign w163 = ~in1[9];
assign w164 = ~in1[9];
assign w165 = ~in1[9];
assign w166 = ~in1[9];
assign w167 = ~in1[9];
assign w168 = ~in1[9];
assign w169 = ~in1[9];
assign w170 = ~in1[9];
assign w171 = ~in1[9];
assign w172 = ~in1[9];
assign w173 = ~in1[9];
assign w174 = ~in1[9];
assign w175 = ~in1[9];
assign w176 = in1[10] ~^ in1[9];
assign w177 = in1[10] ~| in1[9];
assign w178 = ~in1[10];
assign w179 = ~in1[10];
assign w180 = ~in1[10];
assign w181 = ~in1[10];
assign w182 = ~in1[10];
assign w183 = ~in1[10];
assign w184 = ~in1[10];
assign w185 = ~in1[10];
assign w186 = ~in1[10];
assign w187 = ~in1[10];
assign w188 = ~in1[10];
assign w189 = ~in1[10];
assign w190 = ~in1[10];
assign w191 = ~in1[10];
assign w192 = ~in1[10];
assign w193 = ~in1[10];
assign w194 = in1[11] ~^ in1[10];
assign w195 = in1[11] ~| in1[10];
assign w196 = ~in1[11];
assign w197 = ~in1[11];
assign w198 = ~in1[11];
assign w199 = ~in1[11];
assign w200 = ~in1[11];
assign w201 = ~in1[11];
assign w202 = ~in1[11];
assign w203 = ~in1[11];
assign w204 = ~in1[11];
assign w205 = ~in1[11];
assign w206 = ~in1[11];
assign w207 = ~in1[11];
assign w208 = ~in1[11];
assign w209 = ~in1[11];
assign w210 = ~in1[11];
assign w211 = ~in1[11];
assign w212 = in1[12] ~^ in1[11];
assign w213 = in1[12] ~| in1[11];
assign w214 = ~in1[12];
assign w215 = ~in1[12];
assign w216 = ~in1[12];
assign w217 = ~in1[12];
assign w218 = ~in1[12];
assign w219 = ~in1[12];
assign w220 = ~in1[12];
assign w221 = ~in1[12];
assign w222 = ~in1[12];
assign w223 = ~in1[12];
assign w224 = ~in1[12];
assign w225 = ~in1[12];
assign w226 = ~in1[12];
assign w227 = ~in1[12];
assign w228 = ~in1[12];
assign w229 = ~in1[12];
assign w230 = in1[13] ~^ in1[12];
assign w231 = in1[13] ~| in1[12];
assign w232 = ~in1[13];
assign w233 = ~in1[13];
assign w234 = ~in1[13];
assign w235 = ~in1[13];
assign w236 = ~in1[13];
assign w237 = ~in1[13];
assign w238 = ~in1[13];
assign w239 = ~in1[13];
assign w240 = ~in1[13];
assign w241 = ~in1[13];
assign w242 = ~in1[13];
assign w243 = ~in1[13];
assign w244 = ~in1[13];
assign w245 = ~in1[13];
assign w246 = ~in1[13];
assign w247 = ~in1[13];
assign w248 = in1[14] ~^ in1[13];
assign w249 = in1[14] ~| in1[13];
assign w250 = ~in1[14];
assign w251 = ~in1[14];
assign w252 = ~in1[14];
assign w253 = ~in1[14];
assign w254 = ~in1[14];
assign w255 = ~in1[14];
assign w256 = ~in1[14];
assign w257 = ~in1[14];
assign w258 = ~in1[14];
assign w259 = ~in1[14];
assign w260 = ~in1[14];
assign w261 = ~in1[14];
assign w262 = ~in1[14];
assign w263 = ~in1[14];
assign w264 = ~in1[14];
assign w265 = ~in1[14];
assign w266 = in1[15] ~^ in1[14];
assign w267 = in1[15] ~| in1[14];
assign w268 = ~in1[15];
assign w269 = ~in1[15];
assign w270 = ~in1[15];
assign w271 = ~in1[15];
assign w272 = ~in1[15];
assign w273 = ~in1[15];
assign w274 = ~in1[15];
assign w275 = ~in1[15];
assign w276 = ~in1[15];
assign w277 = ~in1[15];
assign w278 = ~in1[15];
assign w279 = ~in1[15];
assign w280 = ~in1[15];
assign w281 = ~in1[15];
assign w282 = ~in1[15];
assign w283 = ~in1[15];
assign w284 = in1[16] ~^ in1[15];
assign w285 = in1[16] ~| in1[15];
assign w286 = ~in1[16];
assign w287 = ~in1[16];
assign w288 = ~in1[16];
assign w289 = ~in1[16];
assign w290 = ~in1[16];
assign w291 = ~in1[16];
assign w292 = ~in1[16];
assign w293 = ~in1[16];
assign w294 = ~in1[16];
assign w295 = ~in1[16];
assign w296 = ~in1[16];
assign w297 = ~in1[16];
assign w298 = ~in1[16];
assign w299 = ~in1[16];
assign w300 = ~in1[16];
assign w301 = ~in1[16];
assign w302 = in1[17] ~^ in1[16];
assign w303 = in1[17] ~| in1[16];
assign w304 = ~in1[17];
assign w305 = ~in1[17];
assign w306 = ~in1[17];
assign w307 = ~in1[17];
assign w308 = ~in1[17];
assign w309 = ~in1[17];
assign w310 = ~in1[17];
assign w311 = ~in1[17];
assign w312 = ~in1[17];
assign w313 = ~in1[17];
assign w314 = ~in1[17];
assign w315 = ~in1[17];
assign w316 = ~in1[17];
assign w317 = ~in1[17];
assign w318 = ~in1[17];
assign w319 = ~in1[17];
assign w320 = in1[18] ~^ in1[17];
assign w321 = in1[18] ~| in1[17];
assign w322 = ~in1[18];
assign w323 = ~in1[18];
assign w324 = ~in1[18];
assign w325 = ~in1[18];
assign w326 = ~in1[18];
assign w327 = ~in1[18];
assign w328 = ~in1[18];
assign w329 = ~in1[18];
assign w330 = ~in1[18];
assign w331 = ~in1[18];
assign w332 = ~in1[18];
assign w333 = ~in1[18];
assign w334 = ~in1[18];
assign w335 = ~in1[18];
assign w336 = ~in1[18];
assign w337 = ~in1[18];
assign w338 = in1[19] ~^ in1[18];
assign w339 = in1[19] ~| in1[18];
assign w340 = ~in1[19];
assign w341 = ~in1[19];
assign w342 = ~in1[19];
assign w343 = ~in1[19];
assign w344 = ~in1[19];
assign w345 = ~in1[19];
assign w346 = ~in1[19];
assign w347 = ~in1[19];
assign w348 = ~in1[19];
assign w349 = ~in1[19];
assign w350 = ~in1[19];
assign w351 = ~in1[19];
assign w352 = ~in1[19];
assign w353 = ~in1[19];
assign w354 = ~in1[19];
assign w355 = ~in1[19];
assign w356 = in1[20] ~^ in1[19];
assign w357 = in1[20] ~| in1[19];
assign w358 = ~in1[20];
assign w359 = ~in1[20];
assign w360 = ~in1[20];
assign w361 = ~in1[20];
assign w362 = ~in1[20];
assign w363 = ~in1[20];
assign w364 = ~in1[20];
assign w365 = ~in1[20];
assign w366 = ~in1[20];
assign w367 = ~in1[20];
assign w368 = ~in1[20];
assign w369 = ~in1[20];
assign w370 = ~in1[20];
assign w371 = ~in1[20];
assign w372 = ~in1[20];
assign w373 = ~in1[20];
assign w374 = in1[21] ~^ in1[20];
assign w375 = in1[21] ~| in1[20];
assign w376 = ~in1[21];
assign w377 = ~in1[21];
assign w378 = ~in1[21];
assign w379 = ~in1[21];
assign w380 = ~in1[21];
assign w381 = ~in1[21];
assign w382 = ~in1[21];
assign w383 = ~in1[21];
assign w384 = ~in1[21];
assign w385 = ~in1[21];
assign w386 = ~in1[21];
assign w387 = ~in1[21];
assign w388 = ~in1[21];
assign w389 = ~in1[21];
assign w390 = ~in1[21];
assign w391 = ~in1[21];
assign w392 = in1[22] ~^ in1[21];
assign w393 = in1[22] ~| in1[21];
assign w394 = ~in1[22];
assign w395 = ~in1[22];
assign w396 = ~in1[22];
assign w397 = ~in1[22];
assign w398 = ~in1[22];
assign w399 = ~in1[22];
assign w400 = ~in1[22];
assign w401 = ~in1[22];
assign w402 = ~in1[22];
assign w403 = ~in1[22];
assign w404 = ~in1[22];
assign w405 = ~in1[22];
assign w406 = ~in1[22];
assign w407 = ~in1[22];
assign w408 = ~in1[22];
assign w409 = ~in1[22];
assign w410 = in1[23] ~^ in1[22];
assign w411 = in1[23] ~| in1[22];
assign w412 = ~in1[23];
assign w413 = ~in1[23];
assign w414 = ~in1[23];
assign w415 = ~in1[23];
assign w416 = ~in1[23];
assign w417 = ~in1[23];
assign w418 = ~in1[23];
assign w419 = ~in1[23];
assign w420 = ~in1[23];
assign w421 = ~in1[23];
assign w422 = ~in1[23];
assign w423 = ~in1[23];
assign w424 = ~in1[23];
assign w425 = ~in1[23];
assign w426 = ~in1[23];
assign w427 = ~in1[23];
assign w428 = in1[24] ~^ in1[23];
assign w429 = in1[24] ~| in1[23];
assign w430 = ~in1[24];
assign w431 = ~in1[24];
assign w432 = ~in1[24];
assign w433 = ~in1[24];
assign w434 = ~in1[24];
assign w435 = ~in1[24];
assign w436 = ~in1[24];
assign w437 = ~in1[24];
assign w438 = ~in1[24];
assign w439 = ~in1[24];
assign w440 = ~in1[24];
assign w441 = ~in1[24];
assign w442 = ~in1[24];
assign w443 = ~in1[24];
assign w444 = ~in1[24];
assign w445 = ~in1[24];
assign w446 = in1[25] ~^ in1[24];
assign w447 = in1[25] ~| in1[24];
assign w448 = ~in1[25];
assign w449 = ~in1[25];
assign w450 = ~in1[25];
assign w451 = ~in1[25];
assign w452 = ~in1[25];
assign w453 = ~in1[25];
assign w454 = ~in1[25];
assign w455 = ~in1[25];
assign w456 = ~in1[25];
assign w457 = ~in1[25];
assign w458 = ~in1[25];
assign w459 = ~in1[25];
assign w460 = ~in1[25];
assign w461 = ~in1[25];
assign w462 = ~in1[25];
assign w463 = in1[26] ~^ in1[25];
assign w464 = in1[26] ~| in1[25];
assign w465 = ~in1[26];
assign w466 = ~in1[26];
assign w467 = ~in1[26];
assign w468 = ~in1[26];
assign w469 = ~in1[26];
assign w470 = ~in1[26];
assign w471 = ~in1[26];
assign w472 = ~in1[26];
assign w473 = ~in1[26];
assign w474 = ~in1[26];
assign w475 = ~in1[26];
assign w476 = ~in1[26];
assign w477 = ~in1[26];
assign w478 = ~in1[26];
assign w479 = in1[27] ~^ in1[26];
assign w480 = in1[27] ~| in1[26];
assign w481 = ~in1[27];
assign w482 = ~in1[27];
assign w483 = ~in1[27];
assign w484 = ~in1[27];
assign w485 = ~in1[27];
assign w486 = ~in1[27];
assign w487 = ~in1[27];
assign w488 = ~in1[27];
assign w489 = ~in1[27];
assign w490 = ~in1[27];
assign w491 = ~in1[27];
assign w492 = ~in1[27];
assign w493 = ~in1[27];
assign w494 = in1[28] ~^ in1[27];
assign w495 = in1[28] ~| in1[27];
assign w496 = ~in1[28];
assign w497 = ~in1[28];
assign w498 = ~in1[28];
assign w499 = ~in1[28];
assign w500 = ~in1[28];
assign w501 = ~in1[28];
assign w502 = ~in1[28];
assign w503 = ~in1[28];
assign w504 = ~in1[28];
assign w505 = ~in1[28];
assign w506 = ~in1[28];
assign w507 = ~in1[28];
assign w508 = in1[29] ~^ in1[28];
assign w509 = in1[29] ~| in1[28];
assign w510 = ~in1[29];
assign w511 = ~in1[29];
assign w512 = ~in1[29];
assign w513 = ~in1[29];
assign w514 = ~in1[29];
assign w515 = ~in1[29];
assign w516 = ~in1[29];
assign w517 = ~in1[29];
assign w518 = ~in1[29];
assign w519 = in1[30] ~^ in1[29];
assign w520 = in1[30] ~| in1[29];
assign w521 = ~in1[30];
assign w522 = ~in1[30];
assign w523 = ~in1[30];
assign w524 = ~in1[30];
assign w525 = ~in1[30];
assign w526 = ~in1[30];
assign w527 = ~in1[30];
assign w528 = ~in1[30];
assign w529 = ~in1[30];
assign w530 = in1[31] ~^ in1[30];
assign w531 = in1[31] ~| in1[30];
assign w532 = ~in1[31];
assign w533 = ~in1[31];
assign w534 = ~in1[31];
assign w535 = ~in1[31];
assign w536 = ~in1[31];
assign w537 = ~in1[31];
assign w538 = ~in1[31];
assign w539 = ~in1[31];
assign w540 = ~in2[4];
assign w541 = ~in2[30];
assign w542 = ~in2[31];
assign w543 = ~in3[0];
assign w544 = in3[2] & in2[0];
assign w545 = in3[2] ~| in2[0];
assign w546 = ~in3[2];
assign w547 = ~in3[3];
assign w548 = ~in3[4];
assign w549 = in3[5] ~^ in2[3];
assign w550 = in3[5] | in2[3];
assign w551 = in3[5] & in2[3];
assign w552 = ~in3[5];
assign w553 = ~in3[6];
assign w554 = ~in3[7];
assign w555 = in3[8] ~^ in2[6];
assign w556 = in3[8] | in2[6];
assign w557 = in3[8] & in2[6];
assign w558 = ~in3[8];
assign w559 = ~in3[9];
assign w560 = ~in3[10];
assign w561 = in3[11] ~^ in2[9];
assign w562 = in3[11] | in2[9];
assign w563 = in3[11] & in2[9];
assign w564 = ~in3[11];
assign w565 = ~in3[12];
assign w566 = ~in3[13];
assign w567 = in3[14] ~^ in2[12];
assign w568 = in3[14] & in2[12];
assign w569 = in3[14] | in2[12];
assign w570 = ~in3[14];
assign w571 = ~in3[15];
assign w572 = ~in3[16];
assign w573 = in3[17] ~^ in2[15];
assign w574 = in3[17] | in2[15];
assign w575 = in3[17] & in2[15];
assign w576 = ~in3[17];
assign w577 = ~in3[18];
assign w578 = ~in3[19];
assign w579 = in3[20] ~^ in2[18];
assign w580 = in3[20] & in2[18];
assign w581 = in3[20] | in2[18];
assign w582 = ~in3[20];
assign w583 = ~in3[21];
assign w584 = ~in3[22];
assign w585 = in3[23] ~^ in2[21];
assign w586 = in3[23] & in2[21];
assign w587 = in3[23] | in2[21];
assign w588 = ~in3[23];
assign w589 = ~in3[24];
assign w590 = ~in3[25];
assign w591 = in3[26] ~^ in2[24];
assign w592 = in3[26] & in2[24];
assign w593 = in3[26] | in2[24];
assign w594 = ~in3[26];
assign w595 = ~in3[27];
assign w596 = ~in3[28];
assign w597 = in3[29] ~^ in2[27];
assign w598 = in3[29] | in2[27];
assign w599 = in3[29] & in2[27];
assign w600 = ~in3[29];
assign w601 = in3[30] ~^ in3[29];
assign w602 = ~in3[30];
assign w603 = ~in3[31];
assign w604 = w14 | w22;
assign w605 = w17 | w39;
assign w606 = w34 | w52;
assign w607 = w57 | w75;
assign w608 = w70 | w93;
assign w609 = w96 | w118;
assign w610 = w106 | w129;
assign w611 = w124 | w142;
assign w612 = w147 | w165;
assign w613 = w160 | w178;
assign w614 = w183 | w201;
assign w615 = w196 | w214;
assign w616 = w219 | w232;
assign w617 = w244 | w255;
assign w618 = w255 | w273;
assign w619 = w273 | w293;
assign w620 = w301 | w319;
assign w621 = w307 | w333;
assign w622 = w325 | w345;
assign w623 = w347 | w363;
assign w624 = w371 | w377;
assign w625 = w389 | w395;
assign w626 = w403 | w416;
assign w627 = w417 | w444;
assign w628 = w436 | w461;
assign w629 = w450 | w467;
assign w630 = w474 | w486;
assign w631 = w484 | w500;
assign w632 = w506 | w510;
assign w633 = w512 | w521;
assign w634 = w526 | w533;
assign w635 = in3[1] & w543;
assign w636 = w546 ~| in3[1];
assign w637 = w546 ~^ in3[1];
assign w638 = w547 ~^ in3[2];
assign w639 = w547 ~| in3[4];
assign w640 = w548 | in3[3];
assign w641 = w548 | in3[5];
assign w642 = in3[5] & w548;
assign w643 = w553 ~^ in3[5];
assign w644 = w553 ~| in3[7];
assign w645 = w554 | in3[6];
assign w646 = in3[8] & w554;
assign w647 = w554 | in3[8];
assign w648 = w559 ~^ in3[8];
assign w649 = w559 ~| in3[10];
assign w650 = w560 | in3[9];
assign w651 = in3[11] & w560;
assign w652 = w560 | in3[11];
assign w653 = w565 ~^ in3[11];
assign w654 = w565 ~| in3[13];
assign w655 = w566 | in3[12];
assign w656 = in3[14] & w566;
assign w657 = w566 | in3[14];
assign w658 = w571 ~^ in3[14];
assign w659 = w571 ~| in3[16];
assign w660 = w572 | in3[15];
assign w661 = w572 | in3[17];
assign w662 = in3[17] & w572;
assign w663 = w577 ~^ in3[17];
assign w664 = w577 ~| in3[19];
assign w665 = w578 | in3[18];
assign w666 = w578 | in3[20];
assign w667 = in3[20] & w578;
assign w668 = w583 ~^ in3[20];
assign w669 = w583 ~| in3[22];
assign w670 = w584 | in3[21];
assign w671 = in3[23] & w584;
assign w672 = w584 | in3[23];
assign w673 = w589 ~^ in3[23];
assign w674 = w589 ~| in3[25];
assign w675 = w590 | in3[24];
assign w676 = w590 | in3[26];
assign w677 = in3[26] & w590;
assign w678 = w595 ~^ in3[26];
assign w679 = w595 | in3[28];
assign w680 = w596 | in3[27];
assign w681 = in3[29] & w596;
assign w682 = w596 | in3[29];
assign w683 = in3[31] | w601;
assign w684 = w602 | in3[31];
assign w685 = w601 | w603;
assign w686 = w603 | in3[30];
assign w687 = w602 | w603;
assign w688 = w604 & w605;
assign w689 = ~w635;
assign w690 = ~w635;
assign w691 = ~w635;
assign w692 = ~w635;
assign w693 = ~w635;
assign w694 = ~w635;
assign w695 = ~w635;
assign w696 = ~w635;
assign w697 = ~w635;
assign w698 = ~w635;
assign w699 = ~w635;
assign w700 = ~w635;
assign w701 = ~w635;
assign w702 = ~w635;
assign w703 = ~w635;
assign w704 = ~w635;
assign w705 = w543 & w636;
assign w706 = in3[0] & w637;
assign w707 = ~w637;
assign w708 = in3[2] & w639;
assign w709 = in3[2] ~| w640;
assign w710 = w547 | w641;
assign w711 = ~w641;
assign w712 = ~w642;
assign w713 = in3[5] & w644;
assign w714 = in3[5] ~| w645;
assign w715 = ~w646;
assign w716 = w553 | w647;
assign w717 = ~w647;
assign w718 = in3[8] & w649;
assign w719 = in3[8] ~| w650;
assign w720 = ~w651;
assign w721 = w559 | w652;
assign w722 = ~w652;
assign w723 = in3[11] & w654;
assign w724 = in3[11] ~| w655;
assign w725 = ~w656;
assign w726 = w565 | w657;
assign w727 = ~w657;
assign w728 = in3[14] & w659;
assign w729 = in3[14] ~| w660;
assign w730 = w571 | w661;
assign w731 = ~w661;
assign w732 = ~w662;
assign w733 = in3[17] & w664;
assign w734 = in3[17] ~| w665;
assign w735 = w577 | w666;
assign w736 = ~w666;
assign w737 = ~w667;
assign w738 = in3[20] & w669;
assign w739 = in3[20] ~| w670;
assign w740 = ~w671;
assign w741 = w583 | w672;
assign w742 = ~w672;
assign w743 = in3[23] & w674;
assign w744 = in3[23] ~| w675;
assign w745 = w589 | w676;
assign w746 = ~w676;
assign w747 = ~w677;
assign w748 = w594 | w679;
assign w749 = in3[26] | w680;
assign w750 = ~w681;
assign w751 = w595 | w682;
assign w752 = ~w682;
assign w753 = w274 ~| w683;
assign w754 = w60 | w683;
assign w755 = w240 | w683;
assign w756 = w204 | w683;
assign w757 = w222 | w683;
assign w758 = w42 | w683;
assign w759 = w258 | w683;
assign w760 = w132 | w683;
assign w761 = w108 ~| w683;
assign w762 = w186 | w683;
assign w763 = w78 | w683;
assign w764 = w25 | w683;
assign w765 = w150 | w683;
assign w766 = w168 | w683;
assign w767 = w101 | w683;
assign w768 = w600 | w684;
assign w769 = w683 & w685;
assign w770 = w16 | w685;
assign w771 = in3[29] | w686;
assign w772 = w600 | w687;
assign w773 = w50 ~^ w688;
assign w774 = w51 | w688;
assign w775 = w300 ~| w689;
assign w776 = w226 ~| w689;
assign w777 = w29 ~| w690;
assign w778 = w172 ~| w690;
assign w779 = w280 ~| w691;
assign w780 = w261 ~| w691;
assign w781 = w459 ~| w692;
assign w782 = w208 ~| w692;
assign w783 = w319 ~| w693;
assign w784 = w46 ~| w693;
assign w785 = w497 ~| w694;
assign w786 = w478 ~| w694;
assign w787 = w102 ~| w695;
assign w788 = w121 ~| w695;
assign w789 = w353 ~| w696;
assign w790 = w387 ~| w696;
assign w791 = w521 ~| w697;
assign w792 = w156 ~| w697;
assign w793 = w493 ~| w698;
assign w794 = w247 ~| w698;
assign w795 = w535 ~| w699;
assign w796 = w138 ~| w699;
assign w797 = w10 ~| w700;
assign w798 = w426 ~| w700;
assign w799 = w372 ~| w701;
assign w800 = w406 ~| w701;
assign w801 = w190 ~| w702;
assign w802 = w82 ~| w702;
assign w803 = w517 ~| w703;
assign w804 = w64 ~| w703;
assign w805 = w335 ~| w704;
assign w806 = w435 ~| w704;
assign w807 = ~w705;
assign w808 = ~w705;
assign w809 = ~w705;
assign w810 = ~w705;
assign w811 = ~w705;
assign w812 = ~w705;
assign w813 = ~w705;
assign w814 = ~w705;
assign w815 = ~w705;
assign w816 = ~w705;
assign w817 = ~w705;
assign w818 = ~w705;
assign w819 = ~w705;
assign w820 = ~w705;
assign w821 = ~w705;
assign w822 = ~w705;
assign w823 = ~w706;
assign w824 = ~w706;
assign w825 = ~w706;
assign w826 = ~w706;
assign w827 = ~w706;
assign w828 = ~w706;
assign w829 = ~w706;
assign w830 = ~w706;
assign w831 = ~w706;
assign w832 = ~w706;
assign w833 = ~w706;
assign w834 = ~w706;
assign w835 = ~w706;
assign w836 = ~w706;
assign w837 = ~w706;
assign w838 = ~w706;
assign w839 = ~w706;
assign w840 = in3[0] & w707;
assign w841 = w708 | w709;
assign w842 = w546 ~| w710;
assign w843 = w642 | w711;
assign w844 = in3[3] ~| w712;
assign w845 = w713 | w714;
assign w846 = in3[6] | w715;
assign w847 = w552 ~| w716;
assign w848 = w646 | w717;
assign w849 = w718 | w719;
assign w850 = in3[9] | w720;
assign w851 = w558 ~| w721;
assign w852 = w651 | w722;
assign w853 = w723 | w724;
assign w854 = in3[12] | w725;
assign w855 = w564 ~| w726;
assign w856 = w656 | w727;
assign w857 = w728 | w729;
assign w858 = w570 ~| w730;
assign w859 = w662 | w731;
assign w860 = in3[15] | w732;
assign w861 = w733 | w734;
assign w862 = w576 ~| w735;
assign w863 = w667 | w736;
assign w864 = in3[18] | w737;
assign w865 = w738 | w739;
assign w866 = in3[21] | w740;
assign w867 = w582 ~| w741;
assign w868 = w671 | w742;
assign w869 = w743 | w744;
assign w870 = w588 ~| w745;
assign w871 = w677 | w746;
assign w872 = in3[24] | w747;
assign w873 = w748 & w749;
assign w874 = in3[27] | w750;
assign w875 = w594 | w751;
assign w876 = w681 | w752;
assign w877 = w6 | w769;
assign w878 = w768 & w771;
assign w879 = w114 | w772;
assign w880 = w201 | w772;
assign w881 = w165 | w772;
assign w882 = w22 | w772;
assign w883 = w101 | w772;
assign w884 = w240 ~| w772;
assign w885 = w219 | w772;
assign w886 = w147 | w772;
assign w887 = w183 | w772;
assign w888 = w129 | w772;
assign w889 = w57 | w772;
assign w890 = w75 | w772;
assign w891 = w9 | w772;
assign w892 = w39 | w772;
assign w893 = w685 ~| w773;
assign w894 = w606 & w774;
assign w895 = w378 ~| w807;
assign w896 = w94 ~| w807;
assign w897 = w274 ~| w808;
assign w898 = w130 ~| w808;
assign w899 = w364 ~| w809;
assign w900 = w58 ~| w809;
assign w901 = w23 ~| w810;
assign w902 = w202 ~| w810;
assign w903 = w400 ~| w811;
assign w904 = w110 ~| w811;
assign w905 = w2 ~| w812;
assign w906 = w290 ~| w812;
assign w907 = w250 ~| w813;
assign w908 = w76 ~| w813;
assign w909 = w432 ~| w814;
assign w910 = w512 ~| w814;
assign w911 = w526 ~| w815;
assign w912 = w327 ~| w815;
assign w913 = w236 ~| w816;
assign w914 = w184 ~| w816;
assign w915 = w498 ~| w817;
assign w916 = w166 ~| w817;
assign w917 = w344 ~| w818;
assign w918 = w534 ~| w818;
assign w919 = w452 ~| w819;
assign w920 = w471 ~| w819;
assign w921 = w148 ~| w820;
assign w922 = w40 ~| w820;
assign w923 = w304 ~| w821;
assign w924 = w220 ~| w821;
assign w925 = w418 ~| w822;
assign w926 = w484 ~| w822;
assign w927 = w773 ~| w832;
assign w928 = w16 ~| w833;
assign w929 = ~w840;
assign w930 = ~w840;
assign w931 = ~w840;
assign w932 = ~w840;
assign w933 = ~w840;
assign w934 = ~w840;
assign w935 = ~w840;
assign w936 = ~w840;
assign w937 = ~w840;
assign w938 = ~w840;
assign w939 = ~w840;
assign w940 = ~w840;
assign w941 = ~w840;
assign w942 = ~w840;
assign w943 = ~w840;
assign w944 = ~w840;
assign w945 = ~w841;
assign w946 = ~w841;
assign w947 = ~w841;
assign w948 = ~w841;
assign w949 = ~w841;
assign w950 = ~w841;
assign w951 = ~w841;
assign w952 = ~w841;
assign w953 = ~w841;
assign w954 = ~w841;
assign w955 = ~w841;
assign w956 = ~w841;
assign w957 = ~w841;
assign w958 = ~w841;
assign w959 = ~w841;
assign w960 = ~w841;
assign w961 = w638 & w843;
assign w962 = ~w843;
assign w963 = w546 & w844;
assign w964 = ~w845;
assign w965 = ~w845;
assign w966 = ~w845;
assign w967 = ~w845;
assign w968 = ~w845;
assign w969 = ~w845;
assign w970 = ~w845;
assign w971 = ~w845;
assign w972 = ~w845;
assign w973 = ~w845;
assign w974 = ~w845;
assign w975 = ~w845;
assign w976 = ~w845;
assign w977 = ~w845;
assign w978 = ~w845;
assign w979 = ~w845;
assign w980 = in3[5] ~| w846;
assign w981 = w643 & w848;
assign w982 = ~w848;
assign w983 = ~w849;
assign w984 = ~w849;
assign w985 = ~w849;
assign w986 = ~w849;
assign w987 = ~w849;
assign w988 = ~w849;
assign w989 = ~w849;
assign w990 = ~w849;
assign w991 = ~w849;
assign w992 = ~w849;
assign w993 = ~w849;
assign w994 = ~w849;
assign w995 = ~w849;
assign w996 = ~w849;
assign w997 = ~w849;
assign w998 = ~w849;
assign w999 = in3[8] ~| w850;
assign w1000 = w648 & w852;
assign w1001 = ~w852;
assign w1002 = ~w853;
assign w1003 = ~w853;
assign w1004 = ~w853;
assign w1005 = ~w853;
assign w1006 = ~w853;
assign w1007 = ~w853;
assign w1008 = ~w853;
assign w1009 = ~w853;
assign w1010 = ~w853;
assign w1011 = ~w853;
assign w1012 = ~w853;
assign w1013 = ~w853;
assign w1014 = ~w853;
assign w1015 = ~w853;
assign w1016 = ~w853;
assign w1017 = ~w853;
assign w1018 = in3[11] ~| w854;
assign w1019 = w653 & w856;
assign w1020 = ~w856;
assign w1021 = ~w857;
assign w1022 = ~w857;
assign w1023 = ~w857;
assign w1024 = ~w857;
assign w1025 = ~w857;
assign w1026 = ~w857;
assign w1027 = ~w857;
assign w1028 = ~w857;
assign w1029 = ~w857;
assign w1030 = ~w857;
assign w1031 = ~w857;
assign w1032 = ~w857;
assign w1033 = ~w857;
assign w1034 = ~w857;
assign w1035 = ~w857;
assign w1036 = ~w857;
assign w1037 = w658 & w859;
assign w1038 = ~w859;
assign w1039 = in3[14] ~| w860;
assign w1040 = ~w861;
assign w1041 = ~w861;
assign w1042 = ~w861;
assign w1043 = ~w861;
assign w1044 = ~w861;
assign w1045 = ~w861;
assign w1046 = ~w861;
assign w1047 = ~w861;
assign w1048 = ~w861;
assign w1049 = ~w861;
assign w1050 = ~w861;
assign w1051 = ~w861;
assign w1052 = w663 & w863;
assign w1053 = ~w863;
assign w1054 = in3[17] ~| w864;
assign w1055 = ~w865;
assign w1056 = ~w865;
assign w1057 = ~w865;
assign w1058 = ~w865;
assign w1059 = ~w865;
assign w1060 = ~w865;
assign w1061 = ~w865;
assign w1062 = ~w865;
assign w1063 = ~w865;
assign w1064 = ~w865;
assign w1065 = ~w865;
assign w1066 = ~w865;
assign w1067 = in3[20] ~| w866;
assign w1068 = w668 & w868;
assign w1069 = ~w868;
assign w1070 = ~w869;
assign w1071 = ~w869;
assign w1072 = ~w869;
assign w1073 = ~w869;
assign w1074 = ~w869;
assign w1075 = ~w869;
assign w1076 = ~w869;
assign w1077 = ~w869;
assign w1078 = ~w869;
assign w1079 = w673 & w871;
assign w1080 = ~w871;
assign w1081 = in3[23] ~| w872;
assign w1082 = w27 ~| w873;
assign w1083 = w264 ~| w873;
assign w1084 = w185 ~| w873;
assign w1085 = w298 ~| w873;
assign w1086 = w97 ~| w873;
assign w1087 = w154 ~| w873;
assign w1088 = w161 ~| w873;
assign w1089 = w112 ~| w873;
assign w1090 = w206 ~| w873;
assign w1091 = w278 ~| w873;
assign w1092 = w35 ~| w873;
assign w1093 = w52 ~| w873;
assign w1094 = w11 ~| w873;
assign w1095 = w136 ~| w873;
assign w1096 = w71 ~| w873;
assign w1097 = w232 ~| w873;
assign w1098 = w316 ~| w873;
assign w1099 = w221 ~| w873;
assign w1100 = in3[26] | w874;
assign w1101 = w678 & w876;
assign w1102 = ~w876;
assign w1103 = w877 ~^ in2[30];
assign w1104 = w541 | w877;
assign w1105 = w41 ~| w878;
assign w1106 = w31 ~| w878;
assign w1107 = w200 ~| w878;
assign w1108 = w1 | w878;
assign w1109 = w133 ~| w878;
assign w1110 = w67 ~| w878;
assign w1111 = w108 ~| w878;
assign w1112 = w238 ~| w878;
assign w1113 = w93 | w878;
assign w1114 = w79 ~| w878;
assign w1115 = w192 ~| w878;
assign w1116 = w259 ~| w878;
assign w1117 = w221 ~| w878;
assign w1118 = w162 ~| w878;
assign w1119 = w149 ~| w878;
assign w1120 = w765 & w879;
assign w1121 = w755 & w880;
assign w1122 = w756 & w881;
assign w1123 = w754 & w882;
assign w1124 = w760 & w883;
assign w1125 = w753 | w884;
assign w1126 = w759 & w885;
assign w1127 = w762 & w886;
assign w1128 = w757 & w887;
assign w1129 = w766 & w888;
assign w1130 = w767 & w889;
assign w1131 = w758 & w891;
assign w1132 = w763 & w892;
assign w1133 = w68 ~^ w894;
assign w1134 = w69 | w894;
assign w1135 = w800 | w895;
assign w1136 = w788 | w896;
assign w1137 = w775 | w897;
assign w1138 = w792 | w898;
assign w1139 = w790 | w899;
assign w1140 = w802 | w900;
assign w1141 = w784 | w901;
assign w1142 = w776 | w902;
assign w1143 = w798 | w903;
assign w1144 = w796 | w904;
assign w1145 = w777 | w905;
assign w1146 = w783 | w906;
assign w1147 = w779 | w907;
assign w1148 = w787 | w908;
assign w1149 = w781 | w909;
assign w1150 = w791 | w910;
assign w1151 = w795 | w911;
assign w1152 = w789 | w912;
assign w1153 = w780 | w913;
assign w1154 = w782 | w914;
assign w1155 = w803 | w915;
assign w1156 = w801 | w916;
assign w1157 = w799 | w917;
assign w1158 = w786 | w919;
assign w1159 = w793 | w920;
assign w1160 = w778 | w921;
assign w1161 = w804 | w922;
assign w1162 = w805 | w923;
assign w1163 = w794 | w924;
assign w1164 = w806 | w925;
assign w1165 = w785 | w926;
assign w1166 = w797 | w928;
assign w1167 = w537 ~| w929;
assign w1168 = w211 ~| w929;
assign w1169 = w30 ~| w930;
assign w1170 = w136 ~| w930;
assign w1171 = w528 ~| w931;
assign w1172 = w142 ~| w931;
assign w1173 = w252 ~| w932;
assign w1174 = w833 & w932;
assign w1175 = w436 ~| w933;
assign w1176 = w234 ~| w933;
assign w1177 = w227 ~| w934;
assign w1178 = w44 ~| w934;
assign w1179 = w313 ~| w935;
assign w1180 = w175 ~| w935;
assign w1181 = w513 ~| w936;
assign w1182 = w501 ~| w936;
assign w1183 = w354 ~| w937;
assign w1184 = w59 ~| w937;
assign w1185 = w288 ~| w938;
assign w1186 = w92 ~| w938;
assign w1187 = w369 ~| w939;
assign w1188 = w120 ~| w939;
assign w1189 = w469 ~| w940;
assign w1190 = w401 ~| w940;
assign w1191 = w333 ~| w941;
assign w1192 = w83 ~| w941;
assign w1193 = w482 ~| w942;
assign w1194 = w382 ~| w942;
assign w1195 = w450 ~| w943;
assign w1196 = w417 ~| w943;
assign w1197 = w277 ~| w944;
assign w1198 = w185 ~| w944;
assign w1199 = w535 ~| w945;
assign w1200 = w154 ~| w945;
assign w1201 = w287 ~| w946;
assign w1202 = w134 ~| w946;
assign w1203 = w523 ~| w947;
assign w1204 = w118 ~| w947;
assign w1205 = w18 ~| w948;
assign w1206 = w77 ~| w948;
assign w1207 = w251 ~| w949;
assign w1208 = w205 ~| w949;
assign w1209 = w486 ~| w950;
assign w1210 = w449 ~| w950;
assign w1211 = w515 ~| w951;
assign w1212 = w169 ~| w951;
assign w1213 = w345 ~| w952;
assign w1214 = w310 ~| w952;
assign w1215 = w376 ~| w953;
assign w1216 = w65 ~| w953;
assign w1217 = w1 ~| w954;
assign w1218 = w427 ~| w954;
assign w1219 = w368 ~| w955;
assign w1220 = w275 ~| w955;
assign w1221 = w327 ~| w956;
assign w1222 = w38 ~| w956;
assign w1223 = w232 ~| w957;
assign w1224 = w95 ~| w957;
assign w1225 = w502 ~| w958;
assign w1226 = w408 ~| w958;
assign w1227 = w466 ~| w959;
assign w1228 = w438 ~| w959;
assign w1229 = w193 ~| w960;
assign w1230 = w215 ~| w960;
assign w1231 = ~w961;
assign w1232 = ~w961;
assign w1233 = ~w961;
assign w1234 = ~w961;
assign w1235 = ~w961;
assign w1236 = ~w961;
assign w1237 = ~w961;
assign w1238 = ~w961;
assign w1239 = ~w961;
assign w1240 = ~w961;
assign w1241 = ~w961;
assign w1242 = ~w961;
assign w1243 = ~w961;
assign w1244 = ~w961;
assign w1245 = ~w961;
assign w1246 = ~w961;
assign w1247 = ~w961;
assign w1248 = w638 & w962;
assign w1249 = w842 | w963;
assign w1250 = w522 ~| w964;
assign w1251 = w84 ~| w964;
assign w1252 = w26 ~| w965;
assign w1253 = w229 ~| w965;
assign w1254 = w539 ~| w966;
assign w1255 = w34 ~| w966;
assign w1256 = w271 ~| w967;
assign w1257 = w62 ~| w967;
assign w1258 = w514 ~| w968;
assign w1259 = w89 ~| w968;
assign w1260 = w328 ~| w969;
assign w1261 = w291 ~| w969;
assign w1262 = w149 ~| w970;
assign w1263 = w131 ~| w970;
assign w1264 = w489 ~| w971;
assign w1265 = w441 ~| w971;
assign w1266 = w372 ~| w972;
assign w1267 = w170 ~| w972;
assign w1268 = w473 ~| w973;
assign w1269 = w407 ~| w973;
assign w1270 = w353 ~| w974;
assign w1271 = w257 ~| w974;
assign w1272 = w305 ~| w975;
assign w1273 = w188 ~| w975;
assign w1274 = w461 ~| w976;
assign w1275 = w422 ~| w976;
assign w1276 = w197 ~| w977;
assign w1277 = w246 ~| w977;
assign w1278 = w4 ~| w978;
assign w1279 = w107 ~| w978;
assign w1280 = w507 ~| w979;
assign w1281 = w380 ~| w979;
assign w1282 = w847 | w980;
assign w1283 = ~w981;
assign w1284 = ~w981;
assign w1285 = ~w981;
assign w1286 = ~w981;
assign w1287 = ~w981;
assign w1288 = ~w981;
assign w1289 = ~w981;
assign w1290 = ~w981;
assign w1291 = ~w981;
assign w1292 = ~w981;
assign w1293 = ~w981;
assign w1294 = ~w981;
assign w1295 = ~w981;
assign w1296 = ~w981;
assign w1297 = ~w981;
assign w1298 = ~w981;
assign w1299 = ~w981;
assign w1300 = w643 & w982;
assign w1301 = w532 ~| w983;
assign w1302 = w228 ~| w983;
assign w1303 = w19 ~| w984;
assign w1304 = w54 ~| w984;
assign w1305 = w524 ~| w985;
assign w1306 = w242 ~| w985;
assign w1307 = w270 ~| w986;
assign w1308 = w146 ~| w986;
assign w1309 = w515 ~| w987;
assign w1310 = w209 ~| w987;
assign w1311 = w335 ~| w988;
assign w1312 = w295 ~| w988;
assign w1313 = w111 ~| w989;
assign w1314 = w80 ~| w989;
assign w1315 = w481 ~| w990;
assign w1316 = w444 ~| w990;
assign w1317 = w360 ~| w991;
assign w1318 = w191 ~| w991;
assign w1319 = w476 ~| w992;
assign w1320 = w404 ~| w992;
assign w1321 = w341 ~| w993;
assign w1322 = w265 ~| w993;
assign w1323 = w309 ~| w994;
assign w1324 = w128 ~| w994;
assign w1325 = w7 ~| w995;
assign w1326 = w164 ~| w995;
assign w1327 = w499 ~| w996;
assign w1328 = w378 ~| w996;
assign w1329 = w455 ~| w997;
assign w1330 = w412 ~| w997;
assign w1331 = w91 ~| w998;
assign w1332 = w43 ~| w998;
assign w1333 = w851 | w999;
assign w1334 = ~w1000;
assign w1335 = ~w1000;
assign w1336 = ~w1000;
assign w1337 = ~w1000;
assign w1338 = ~w1000;
assign w1339 = ~w1000;
assign w1340 = ~w1000;
assign w1341 = ~w1000;
assign w1342 = ~w1000;
assign w1343 = ~w1000;
assign w1344 = ~w1000;
assign w1345 = ~w1000;
assign w1346 = ~w1000;
assign w1347 = ~w1000;
assign w1348 = ~w1000;
assign w1349 = ~w1000;
assign w1350 = ~w1000;
assign w1351 = w648 & w1001;
assign w1352 = w525 ~| w1002;
assign w1353 = w196 ~| w1002;
assign w1354 = w279 ~| w1003;
assign w1355 = w56 ~| w1003;
assign w1356 = w538 ~| w1004;
assign w1357 = w214 ~| w1004;
assign w1358 = w32 ~| w1005;
assign w1359 = w90 ~| w1005;
assign w1360 = w511 ~| w1006;
assign w1361 = w152 ~| w1006;
assign w1362 = w331 ~| w1007;
assign w1363 = w298 ~| w1007;
assign w1364 = w85 ~| w1008;
assign w1365 = w174 ~| w1008;
assign w1366 = w488 ~| w1009;
assign w1367 = w442 ~| w1009;
assign w1368 = w362 ~| w1010;
assign w1369 = w116 ~| w1010;
assign w1370 = w477 ~| w1011;
assign w1371 = w398 ~| w1011;
assign w1372 = w9 ~| w1012;
assign w1373 = w258 ~| w1012;
assign w1374 = w306 ~| w1013;
assign w1375 = w178 ~| w1013;
assign w1376 = w458 ~| w1014;
assign w1377 = w415 ~| w1014;
assign w1378 = w125 ~| w1015;
assign w1379 = w36 ~| w1015;
assign w1380 = w349 ~| w1016;
assign w1381 = w241 ~| w1016;
assign w1382 = w505 ~| w1017;
assign w1383 = w386 ~| w1017;
assign w1384 = w855 | w1018;
assign w1385 = ~w1019;
assign w1386 = ~w1019;
assign w1387 = ~w1019;
assign w1388 = ~w1019;
assign w1389 = ~w1019;
assign w1390 = ~w1019;
assign w1391 = ~w1019;
assign w1392 = ~w1019;
assign w1393 = ~w1019;
assign w1394 = ~w1019;
assign w1395 = ~w1019;
assign w1396 = ~w1019;
assign w1397 = ~w1019;
assign w1398 = ~w1019;
assign w1399 = ~w1019;
assign w1400 = ~w1019;
assign w1401 = ~w1019;
assign w1402 = w653 & w1020;
assign w1403 = w24 ~| w1021;
assign w1404 = w216 ~| w1021;
assign w1405 = w282 ~| w1022;
assign w1406 = w167 ~| w1022;
assign w1407 = w309 ~| w1023;
assign w1408 = w203 ~| w1023;
assign w1409 = w402 ~| w1024;
assign w1410 = w385 ~| w1024;
assign w1411 = w430 ~| w1025;
assign w1412 = w359 ~| w1025;
assign w1413 = w3 ~| w1026;
assign w1414 = w336 ~| w1026;
assign w1415 = w103 ~| w1027;
assign w1416 = w41 ~| w1027;
assign w1417 = w491 ~| w1028;
assign w1418 = w351 ~| w1028;
assign w1419 = w496 ~| w1029;
assign w1420 = w256 ~| w1029;
assign w1421 = w244 ~| w1030;
assign w1422 = w187 ~| w1031;
assign w1423 = w70 ~| w1031;
assign w1424 = w119 ~| w1032;
assign w1425 = w518 ~| w1033;
assign w1426 = w424 ~| w1033;
assign w1427 = w296 ~| w1034;
assign w1428 = w61 ~| w1034;
assign w1429 = w151 ~| w1035;
assign w1430 = w124 ~| w1035;
assign w1431 = w467 ~| w1036;
assign w1432 = w460 ~| w1036;
assign w1433 = ~w1037;
assign w1434 = ~w1037;
assign w1435 = ~w1037;
assign w1436 = ~w1037;
assign w1437 = ~w1037;
assign w1438 = ~w1037;
assign w1439 = ~w1037;
assign w1440 = ~w1037;
assign w1441 = ~w1037;
assign w1442 = ~w1037;
assign w1443 = ~w1037;
assign w1444 = ~w1037;
assign w1445 = ~w1037;
assign w1446 = ~w1037;
assign w1447 = ~w1037;
assign w1448 = w658 & w1038;
assign w1449 = w858 | w1039;
assign w1450 = w160 ~| w1040;
assign w1451 = w454 ~| w1040;
assign w1452 = w24 ~| w1040;
assign w1453 = w260 ~| w1041;
assign w1454 = w269 ~| w1041;
assign w1455 = w198 ~| w1041;
assign w1456 = w233 ~| w1042;
assign w1457 = w419 ~| w1042;
assign w1458 = w182 ~| w1042;
assign w1459 = w131 ~| w1043;
assign w1460 = w224 ~| w1043;
assign w1461 = w292 ~| w1044;
assign w1462 = w115 ~| w1044;
assign w1463 = w474 ~| w1045;
assign w1464 = w388 ~| w1045;
assign w1465 = w396 ~| w1046;
assign w1466 = w370 ~| w1046;
assign w1467 = w317 ~| w1047;
assign w1468 = w59 ~| w1047;
assign w1469 = w342 ~| w1048;
assign w1470 = w12 ~| w1048;
assign w1471 = w157 ~| w1049;
assign w1472 = w98 ~| w1049;
assign w1473 = w323 ~| w1050;
assign w1474 = w72 ~| w1050;
assign w1475 = w434 ~| w1051;
assign w1476 = w49 ~| w1051;
assign w1477 = ~w1052;
assign w1478 = ~w1052;
assign w1479 = ~w1052;
assign w1480 = ~w1052;
assign w1481 = ~w1052;
assign w1482 = ~w1052;
assign w1483 = ~w1052;
assign w1484 = ~w1052;
assign w1485 = ~w1052;
assign w1486 = ~w1052;
assign w1487 = ~w1052;
assign w1488 = ~w1052;
assign w1489 = ~w1052;
assign w1490 = ~w1052;
assign w1491 = w663 & w1053;
assign w1492 = w862 | w1054;
assign w1493 = w394 ~| w1055;
assign w1494 = w281 ~| w1055;
assign w1495 = w297 ~| w1056;
assign w1496 = w77 ~| w1056;
assign w1497 = w100 ~| w1057;
assign w1498 = w167 ~| w1057;
assign w1499 = w367 ~| w1058;
assign w1500 = w218 ~| w1058;
assign w1501 = w314 ~| w1059;
assign w1502 = w47 ~| w1059;
assign w1503 = w390 ~| w1060;
assign w1504 = w126 ~| w1060;
assign w1505 = w346 ~| w1061;
assign w1506 = w262 ~| w1061;
assign w1507 = w144 ~| w1062;
assign w1508 = w180 ~| w1062;
assign w1509 = w13 ~| w1063;
assign w1510 = w17 ~| w1063;
assign w1511 = w421 ~| w1064;
assign w1512 = w332 ~| w1064;
assign w1513 = w203 ~| w1065;
assign w1514 = w66 ~| w1065;
assign w1515 = w237 ~| w1066;
assign w1516 = w106 ~| w1066;
assign w1517 = w867 | w1067;
assign w1518 = ~w1068;
assign w1519 = ~w1068;
assign w1520 = ~w1068;
assign w1521 = ~w1068;
assign w1522 = ~w1068;
assign w1523 = ~w1068;
assign w1524 = ~w1068;
assign w1525 = ~w1068;
assign w1526 = ~w1068;
assign w1527 = ~w1068;
assign w1528 = ~w1068;
assign w1529 = ~w1068;
assign w1530 = w668 & w1069;
assign w1531 = w15 ~| w1070;
assign w1532 = w289 ~| w1070;
assign w1533 = w21 ~| w1071;
assign w1534 = w350 ~| w1071;
assign w1535 = w272 ~| w1072;
assign w1536 = w48 ~| w1072;
assign w1537 = w143 ~| w1073;
assign w1538 = w113 ~| w1073;
assign w1539 = w210 ~| w1074;
assign w1540 = w245 ~| w1074;
assign w1541 = w223 ~| w1074;
assign w1542 = w324 ~| w1075;
assign w1543 = w318 ~| w1075;
assign w1544 = w74 ~| w1075;
assign w1545 = w139 ~| w1076;
assign w1546 = w53 ~| w1076;
assign w1547 = w95 ~| w1076;
assign w1548 = w364 ~| w1077;
assign w1549 = w179 ~| w1077;
assign w1550 = w254 ~| w1078;
assign w1551 = w173 ~| w1078;
assign w1552 = ~w1079;
assign w1553 = ~w1079;
assign w1554 = ~w1079;
assign w1555 = ~w1079;
assign w1556 = ~w1079;
assign w1557 = ~w1079;
assign w1558 = ~w1079;
assign w1559 = ~w1079;
assign w1560 = ~w1079;
assign w1561 = ~w1079;
assign w1562 = w673 & w1080;
assign w1563 = w870 | w1081;
assign w1564 = w875 & w1100;
assign w1565 = ~w1101;
assign w1566 = ~w1101;
assign w1567 = ~w1101;
assign w1568 = ~w1101;
assign w1569 = ~w1101;
assign w1570 = ~w1101;
assign w1571 = ~w1101;
assign w1572 = ~w1101;
assign w1573 = w678 & w1102;
assign w1574 = w1104 ~^ in2[31];
assign w1575 = w893 ~| w1105;
assign w1576 = w764 & w1108;
assign w1577 = w890 & w1113;
assign w1578 = w839 ~| w1133;
assign w1579 = w685 ~| w1133;
assign w1580 = w607 & w1134;
assign w1581 = w1166 | w1169;
assign w1582 = w8 | w1174;
assign w1583 = w927 | w1184;
assign w1584 = w773 ~| w1240;
assign w1585 = w16 ~| w1241;
assign w1586 = w1133 ~| w1247;
assign w1587 = ~w1248;
assign w1588 = ~w1248;
assign w1589 = ~w1248;
assign w1590 = ~w1248;
assign w1591 = ~w1248;
assign w1592 = ~w1248;
assign w1593 = ~w1248;
assign w1594 = ~w1248;
assign w1595 = ~w1248;
assign w1596 = ~w1248;
assign w1597 = ~w1248;
assign w1598 = ~w1248;
assign w1599 = ~w1248;
assign w1600 = ~w1248;
assign w1601 = ~w1248;
assign w1602 = ~w1248;
assign w1603 = ~w1249;
assign w1604 = ~w1249;
assign w1605 = ~w1249;
assign w1606 = ~w1249;
assign w1607 = ~w1249;
assign w1608 = ~w1249;
assign w1609 = ~w1249;
assign w1610 = ~w1249;
assign w1611 = ~w1249;
assign w1612 = ~w1249;
assign w1613 = ~w1249;
assign w1614 = ~w1249;
assign w1615 = ~w1249;
assign w1616 = ~w1249;
assign w1617 = ~w1249;
assign w1618 = ~w1249;
assign w1619 = ~w1282;
assign w1620 = ~w1282;
assign w1621 = ~w1282;
assign w1622 = ~w1282;
assign w1623 = ~w1282;
assign w1624 = ~w1282;
assign w1625 = ~w1282;
assign w1626 = ~w1282;
assign w1627 = ~w1282;
assign w1628 = ~w1282;
assign w1629 = ~w1282;
assign w1630 = ~w1282;
assign w1631 = ~w1282;
assign w1632 = ~w1282;
assign w1633 = ~w1282;
assign w1634 = ~w1282;
assign w1635 = w773 ~| w1292;
assign w1636 = w16 ~| w1293;
assign w1637 = w1133 ~| w1299;
assign w1638 = ~w1300;
assign w1639 = ~w1300;
assign w1640 = ~w1300;
assign w1641 = ~w1300;
assign w1642 = ~w1300;
assign w1643 = ~w1300;
assign w1644 = ~w1300;
assign w1645 = ~w1300;
assign w1646 = ~w1300;
assign w1647 = ~w1300;
assign w1648 = ~w1300;
assign w1649 = ~w1300;
assign w1650 = ~w1300;
assign w1651 = ~w1300;
assign w1652 = ~w1300;
assign w1653 = ~w1300;
assign w1654 = ~w1333;
assign w1655 = ~w1333;
assign w1656 = ~w1333;
assign w1657 = ~w1333;
assign w1658 = ~w1333;
assign w1659 = ~w1333;
assign w1660 = ~w1333;
assign w1661 = ~w1333;
assign w1662 = ~w1333;
assign w1663 = ~w1333;
assign w1664 = ~w1333;
assign w1665 = ~w1333;
assign w1666 = ~w1333;
assign w1667 = ~w1333;
assign w1668 = ~w1333;
assign w1669 = ~w1333;
assign w1670 = w773 ~| w1343;
assign w1671 = w16 ~| w1344;
assign w1672 = w1133 ~| w1350;
assign w1673 = ~w1351;
assign w1674 = ~w1351;
assign w1675 = ~w1351;
assign w1676 = ~w1351;
assign w1677 = ~w1351;
assign w1678 = ~w1351;
assign w1679 = ~w1351;
assign w1680 = ~w1351;
assign w1681 = ~w1351;
assign w1682 = ~w1351;
assign w1683 = ~w1351;
assign w1684 = ~w1351;
assign w1685 = ~w1351;
assign w1686 = ~w1351;
assign w1687 = ~w1351;
assign w1688 = ~w1351;
assign w1689 = ~w1384;
assign w1690 = ~w1384;
assign w1691 = ~w1384;
assign w1692 = ~w1384;
assign w1693 = ~w1384;
assign w1694 = ~w1384;
assign w1695 = ~w1384;
assign w1696 = ~w1384;
assign w1697 = ~w1384;
assign w1698 = ~w1384;
assign w1699 = ~w1384;
assign w1700 = ~w1384;
assign w1701 = ~w1384;
assign w1702 = ~w1384;
assign w1703 = ~w1384;
assign w1704 = ~w1384;
assign w1705 = w773 ~| w1394;
assign w1706 = w16 ~| w1395;
assign w1707 = w1133 ~| w1401;
assign w1708 = ~w1402;
assign w1709 = ~w1402;
assign w1710 = ~w1402;
assign w1711 = ~w1402;
assign w1712 = ~w1402;
assign w1713 = ~w1402;
assign w1714 = ~w1402;
assign w1715 = ~w1402;
assign w1716 = ~w1402;
assign w1717 = ~w1402;
assign w1718 = ~w1402;
assign w1719 = ~w1402;
assign w1720 = ~w1402;
assign w1721 = ~w1402;
assign w1722 = ~w1402;
assign w1723 = ~w1402;
assign w1724 = w773 ~| w1433;
assign w1725 = w16 ~| w1437;
assign w1726 = w1133 ~| w1447;
assign w1727 = ~w1448;
assign w1728 = ~w1448;
assign w1729 = ~w1448;
assign w1730 = ~w1448;
assign w1731 = ~w1448;
assign w1732 = ~w1448;
assign w1733 = ~w1448;
assign w1734 = ~w1448;
assign w1735 = ~w1448;
assign w1736 = ~w1448;
assign w1737 = ~w1448;
assign w1738 = ~w1448;
assign w1739 = ~w1448;
assign w1740 = ~w1448;
assign w1741 = ~w1448;
assign w1742 = ~w1448;
assign w1743 = ~w1449;
assign w1744 = ~w1449;
assign w1745 = ~w1449;
assign w1746 = ~w1449;
assign w1747 = ~w1449;
assign w1748 = ~w1449;
assign w1749 = ~w1449;
assign w1750 = ~w1449;
assign w1751 = ~w1449;
assign w1752 = ~w1449;
assign w1753 = ~w1449;
assign w1754 = ~w1449;
assign w1755 = ~w1449;
assign w1756 = ~w1449;
assign w1757 = ~w1449;
assign w1758 = w16 ~| w1480;
assign w1759 = w773 ~| w1483;
assign w1760 = w1133 ~| w1489;
assign w1761 = ~w1491;
assign w1762 = ~w1491;
assign w1763 = ~w1491;
assign w1764 = ~w1491;
assign w1765 = ~w1491;
assign w1766 = ~w1491;
assign w1767 = ~w1491;
assign w1768 = ~w1491;
assign w1769 = ~w1491;
assign w1770 = ~w1491;
assign w1771 = ~w1491;
assign w1772 = ~w1491;
assign w1773 = ~w1491;
assign w1774 = ~w1491;
assign w1775 = ~w1492;
assign w1776 = ~w1492;
assign w1777 = ~w1492;
assign w1778 = ~w1492;
assign w1779 = ~w1492;
assign w1780 = ~w1492;
assign w1781 = ~w1492;
assign w1782 = ~w1492;
assign w1783 = ~w1492;
assign w1784 = ~w1492;
assign w1785 = ~w1492;
assign w1786 = ~w1492;
assign w1787 = ~w1492;
assign w1788 = ~w1492;
assign w1789 = ~w1517;
assign w1790 = ~w1517;
assign w1791 = ~w1517;
assign w1792 = ~w1517;
assign w1793 = ~w1517;
assign w1794 = ~w1517;
assign w1795 = ~w1517;
assign w1796 = ~w1517;
assign w1797 = ~w1517;
assign w1798 = ~w1517;
assign w1799 = ~w1517;
assign w1800 = ~w1517;
assign w1801 = w773 ~| w1525;
assign w1802 = w16 ~| w1526;
assign w1803 = w1133 ~| w1528;
assign w1804 = ~w1530;
assign w1805 = ~w1530;
assign w1806 = ~w1530;
assign w1807 = ~w1530;
assign w1808 = ~w1530;
assign w1809 = ~w1530;
assign w1810 = ~w1530;
assign w1811 = ~w1530;
assign w1812 = ~w1530;
assign w1813 = ~w1530;
assign w1814 = ~w1530;
assign w1815 = ~w1530;
assign w1816 = w773 ~| w1554;
assign w1817 = w1133 ~| w1556;
assign w1818 = w16 ~| w1559;
assign w1819 = ~w1562;
assign w1820 = ~w1562;
assign w1821 = ~w1562;
assign w1822 = ~w1562;
assign w1823 = ~w1562;
assign w1824 = ~w1562;
assign w1825 = ~w1562;
assign w1826 = ~w1562;
assign w1827 = ~w1562;
assign w1828 = ~w1562;
assign w1829 = ~w1563;
assign w1830 = ~w1563;
assign w1831 = ~w1563;
assign w1832 = ~w1563;
assign w1833 = ~w1563;
assign w1834 = ~w1563;
assign w1835 = ~w1563;
assign w1836 = ~w1563;
assign w1837 = w128 ~| w1564;
assign w1838 = w256 ~| w1564;
assign w1839 = w107 ~| w1564;
assign w1840 = w204 ~| w1564;
assign w1841 = w233 ~| w1564;
assign w1842 = w180 ~| w1564;
assign w1843 = w81 ~| w1564;
assign w1844 = w45 ~| w1564;
assign w1845 = w223 ~| w1564;
assign w1846 = w88 ~| w1564;
assign w1847 = w168 ~| w1564;
assign w1848 = w18 ~| w1564;
assign w1849 = w143 ~| w1564;
assign w1850 = w287 ~| w1564;
assign w1851 = w271 ~| w1564;
assign w1852 = w10 ~| w1564;
assign w1853 = w55 ~| w1564;
assign w1854 = w773 ~| w1566;
assign w1855 = w1133 ~| w1570;
assign w1856 = w16 ~| w1571;
assign w1857 = ~w1573;
assign w1858 = ~w1573;
assign w1859 = ~w1573;
assign w1860 = ~w1573;
assign w1861 = ~w1573;
assign w1862 = ~w1573;
assign w1863 = ~w1573;
assign w1864 = ~w1573;
assign w1865 = w1123 & w1575;
assign w1866 = w770 & w1576;
assign w1867 = w1192 | w1578;
assign w1868 = w1110 ~| w1579;
assign w1869 = w86 ~^ w1580;
assign w1870 = w87 | w1580;
assign w1871 = w546 ~^ w1581;
assign w1872 = w546 ~^ w1582;
assign w1873 = w1141 ~| w1583;
assign w1874 = w1217 | w1585;
assign w1875 = w533 ~| w1587;
assign w1876 = w39 ~| w1587;
assign w1877 = w283 ~| w1588;
assign w1878 = w165 ~| w1588;
assign w1879 = w523 ~| w1589;
assign w1880 = w129 ~| w1589;
assign w1881 = w261 ~| w1590;
assign w1882 = w1241 & w1590;
assign w1883 = w439 ~| w1591;
assign w1884 = w247 ~| w1591;
assign w1885 = w93 ~| w1592;
assign w1886 = w112 ~| w1592;
assign w1887 = w311 ~| w1593;
assign w1888 = w183 ~| w1593;
assign w1889 = w511 ~| w1594;
assign w1890 = w500 ~| w1594;
assign w1891 = w348 ~| w1595;
assign w1892 = w147 ~| w1595;
assign w1893 = w286 ~| w1596;
assign w1894 = w75 ~| w1596;
assign w1895 = w366 ~| w1597;
assign w1896 = w219 ~| w1597;
assign w1897 = w476 ~| w1598;
assign w1898 = w399 ~| w1598;
assign w1899 = w330 ~| w1599;
assign w1900 = w57 ~| w1599;
assign w1901 = w481 ~| w1600;
assign w1902 = w377 ~| w1600;
assign w1903 = w462 ~| w1601;
assign w1904 = w418 ~| w1601;
assign w1905 = w28 ~| w1602;
assign w1906 = w201 ~| w1602;
assign w1907 = w532 ~| w1603;
assign w1908 = w182 ~| w1603;
assign w1909 = w268 ~| w1604;
assign w1910 = w67 ~| w1604;
assign w1911 = w525 ~| w1605;
assign w1912 = w218 ~| w1605;
assign w1913 = w21 ~| w1606;
assign w1914 = w89 ~| w1606;
assign w1915 = w516 ~| w1607;
assign w1916 = w72 ~| w1607;
assign w1917 = w322 ~| w1608;
assign w1918 = w289 ~| w1608;
assign w1919 = w162 ~| w1609;
assign w1920 = w205 ~| w1609;
assign w1921 = w492 ~| w1610;
assign w1922 = w438 ~| w1610;
assign w1923 = w341 ~| w1611;
assign w1924 = w265 ~| w1611;
assign w1925 = w315 ~| w1612;
assign w1926 = w35 ~| w1612;
assign w1927 = w366 ~| w1613;
assign w1928 = w237 ~| w1613;
assign w1929 = w470 ~| w1614;
assign w1930 = w395 ~| w1614;
assign w1931 = w12 ~| w1615;
assign w1932 = w132 ~| w1615;
assign w1933 = w505 ~| w1616;
assign w1934 = w380 ~| w1616;
assign w1935 = w453 ~| w1617;
assign w1936 = w412 ~| w1617;
assign w1937 = w151 ~| w1618;
assign w1938 = w119 ~| w1618;
assign w1939 = w537 ~| w1619;
assign w1940 = w61 ~| w1619;
assign w1941 = w25 ~| w1620;
assign w1942 = w179 ~| w1620;
assign w1943 = w529 ~| w1621;
assign w1944 = w79 ~| w1621;
assign w1945 = w269 ~| w1622;
assign w1946 = w234 ~| w1622;
assign w1947 = w367 ~| w1623;
assign w1948 = w126 ~| w1623;
assign w1949 = w330 ~| w1624;
assign w1950 = w286 ~| w1624;
assign w1951 = w37 ~| w1625;
assign w1952 = w211 ~| w1625;
assign w1953 = w497 ~| w1626;
assign w1954 = w455 ~| w1626;
assign w1955 = w8 ~| w1627;
assign w1956 = w260 ~| w1627;
assign w1957 = w308 ~| w1628;
assign w1958 = w92 ~| w1628;
assign w1959 = w382 ~| w1629;
assign w1960 = w161 ~| w1629;
assign w1961 = w482 ~| w1630;
assign w1962 = w422 ~| w1630;
assign w1963 = w470 ~| w1631;
assign w1964 = w440 ~| w1631;
assign w1965 = w225 ~| w1632;
assign w1966 = w111 ~| w1632;
assign w1967 = w342 ~| w1633;
assign w1968 = w150 ~| w1633;
assign w1969 = w510 ~| w1634;
assign w1970 = w402 ~| w1634;
assign w1971 = w1278 | w1636;
assign w1972 = w538 ~| w1638;
assign w1973 = w135 ~| w1638;
assign w1974 = w301 ~| w1639;
assign w1975 = w99 ~| w1639;
assign w1976 = w521 ~| w1640;
assign w1977 = w171 ~| w1640;
assign w1978 = w257 ~| w1641;
assign w1979 = w1293 & w1641;
assign w1980 = w343 ~| w1642;
assign w1981 = w190 ~| w1642;
assign w1982 = w517 ~| w1643;
assign w1983 = w504 ~| w1643;
assign w1984 = w433 ~| w1644;
assign w1985 = w199 ~| w1644;
assign w1986 = w217 ~| w1645;
assign w1987 = w81 ~| w1645;
assign w1988 = w270 ~| w1646;
assign w1989 = w46 ~| w1646;
assign w1990 = w325 ~| w1647;
assign w1991 = w109 ~| w1647;
assign w1992 = w383 ~| w1648;
assign w1993 = w153 ~| w1648;
assign w1994 = w475 ~| w1649;
assign w1995 = w23 ~| w1649;
assign w1996 = w363 ~| w1650;
assign w1997 = w235 ~| w1650;
assign w1998 = w488 ~| w1651;
assign w1999 = w404 ~| w1651;
assign w2000 = w453 ~| w1652;
assign w2001 = w420 ~| w1652;
assign w2002 = w307 ~| w1653;
assign w2003 = w55 ~| w1653;
assign w2004 = w539 ~| w1654;
assign w2005 = w216 ~| w1654;
assign w2006 = w19 ~| w1655;
assign w2007 = w243 ~| w1655;
assign w2008 = w359 ~| w1656;
assign w2009 = w97 ~| w1656;
assign w2010 = w292 ~| w1657;
assign w2011 = w49 ~| w1657;
assign w2012 = w522 ~| w1658;
assign w2013 = w127 ~| w1658;
assign w2014 = w354 ~| w1659;
assign w2015 = w305 ~| w1659;
assign w2016 = w253 ~| w1660;
assign w2017 = w114 ~| w1660;
assign w2018 = w503 ~| w1661;
assign w2019 = w448 ~| w1661;
assign w2020 = w181 ~| w1662;
assign w2021 = w279 ~| w1662;
assign w2022 = w334 ~| w1663;
assign w2023 = w60 ~| w1663;
assign w2024 = w388 ~| w1664;
assign w2025 = w198 ~| w1664;
assign w2026 = w483 ~| w1665;
assign w2027 = w423 ~| w1665;
assign w2028 = w2 ~| w1666;
assign w2029 = w153 ~| w1666;
assign w2030 = w513 ~| w1667;
assign w2031 = w394 ~| w1667;
assign w2032 = w465 ~| w1668;
assign w2033 = w432 ~| w1668;
assign w2034 = w171 ~| w1669;
assign w2035 = w73 ~| w1669;
assign w2036 = w1325 | w1671;
assign w2037 = w536 ~| w1673;
assign w2038 = w155 ~| w1673;
assign w2039 = w293 ~| w1674;
assign w2040 = w207 ~| w1674;
assign w2041 = w524 ~| w1675;
assign w2042 = w45 ~| w1675;
assign w2043 = w253 ~| w1676;
assign w2044 = w1344 & w1676;
assign w2045 = w347 ~| w1677;
assign w2046 = w64 ~| w1677;
assign w2047 = w512 ~| w1678;
assign w2048 = w503 ~| w1678;
assign w2049 = w443 ~| w1679;
assign w2050 = w73 ~| w1679;
assign w2051 = w243 ~| w1680;
assign w2052 = w117 ~| w1680;
assign w2053 = w390 ~| w1681;
assign w2054 = w137 ~| w1681;
assign w2055 = w337 ~| w1682;
assign w2056 = w163 ~| w1682;
assign w2057 = w282 ~| w1683;
assign w2058 = w189 ~| w1683;
assign w2059 = w472 ~| w1684;
assign w2060 = w27 ~| w1684;
assign w2061 = w451 ~| w1685;
assign w2062 = w425 ~| w1685;
assign w2063 = w312 ~| w1686;
assign w2064 = w101 ~| w1686;
assign w2065 = w361 ~| w1687;
assign w2066 = w226 ~| w1687;
assign w2067 = w492 ~| w1688;
assign w2068 = w409 ~| w1688;
assign w2069 = w529 ~| w1689;
assign w2070 = w83 ~| w1689;
assign w2071 = w251 ~| w1690;
assign w2072 = w360 ~| w1690;
assign w2073 = w534 ~| w1691;
assign w2074 = w191 ~| w1691;
assign w2075 = w281 ~| w1692;
assign w2076 = w56 ~| w1692;
assign w2077 = w199 ~| w1693;
assign w2078 = w120 ~| w1693;
assign w2079 = w489 ~| w1694;
assign w2080 = w434 ~| w1694;
assign w2081 = w510 ~| w1695;
assign w2082 = w246 ~| w1695;
assign w2083 = w306 ~| w1696;
assign w2084 = w32 ~| w1696;
assign w2085 = w348 ~| w1697;
assign w2086 = w43 ~| w1697;
assign w2087 = w477 ~| w1698;
assign w2088 = w408 ~| w1698;
assign w2089 = w6 ~| w1699;
assign w2090 = w163 ~| w1699;
assign w2091 = w299 ~| w1700;
assign w2092 = w227 ~| w1700;
assign w2093 = w448 ~| w1701;
assign w2094 = w414 ~| w1701;
assign w2095 = w145 ~| w1702;
assign w2096 = w135 ~| w1702;
assign w2097 = w323 ~| w1703;
assign w2098 = w96 ~| w1703;
assign w2099 = w496 ~| w1704;
assign w2100 = w384 ~| w1704;
assign w2101 = w1372 | w1706;
assign w2102 = w536 ~| w1708;
assign w2103 = w127 ~| w1708;
assign w2104 = w276 ~| w1709;
assign w2105 = w63 ~| w1709;
assign w2106 = w527 ~| w1710;
assign w2107 = w239 ~| w1710;
assign w2108 = w263 ~| w1711;
assign w2109 = w1395 & w1711;
assign w2110 = w440 ~| w1712;
assign w2111 = w181 ~| w1712;
assign w2112 = w145 ~| w1713;
assign w2113 = w172 ~| w1713;
assign w2114 = w329 ~| w1714;
assign w2115 = w208 ~| w1714;
assign w2116 = w514 ~| w1715;
assign w2117 = w506 ~| w1715;
assign w2118 = w371 ~| w1716;
assign w2119 = w225 ~| w1716;
assign w2120 = w468 ~| w1717;
assign w2121 = w403 ~| w1717;
assign w2122 = w349 ~| w1718;
assign w2123 = w82 ~| w1718;
assign w2124 = w315 ~| w1719;
assign w2125 = w88 ~| w1719;
assign w2126 = w456 ~| w1720;
assign w2127 = w413 ~| w1720;
assign w2128 = w294 ~| w1721;
assign w2129 = w121 ~| w1721;
assign w2130 = w25 ~| w1722;
assign w2131 = w37 ~| w1722;
assign w2132 = w485 ~| w1723;
assign w2133 = w385 ~| w1723;
assign w2134 = w1413 | w1725;
assign w2135 = w491 ~| w1727;
assign w2136 = w96 ~| w1727;
assign w2137 = w275 ~| w1728;
assign w2138 = w1437 & w1728;
assign w2139 = w518 ~| w1729;
assign w2140 = w186 ~| w1729;
assign w2141 = w78 ~| w1730;
assign w2142 = w340 ~| w1731;
assign w2143 = w42 ~| w1731;
assign w2144 = w60 ~| w1732;
assign w2145 = w168 ~| w1732;
assign w2146 = w528 ~| w1733;
assign w2147 = w132 ~| w1733;
assign w2148 = w250 ~| w1734;
assign w2149 = w222 ~| w1734;
assign w2150 = w20 ~| w1735;
assign w2151 = w204 ~| w1735;
assign w2152 = w452 ~| w1736;
assign w2153 = w405 ~| w1736;
assign w2154 = w502 ~| w1737;
assign w2155 = w469 ~| w1737;
assign w2156 = w322 ~| w1738;
assign w2157 = w299 ~| w1738;
assign w2158 = w431 ~| w1739;
assign w2159 = w389 ~| w1739;
assign w2160 = w312 ~| w1740;
assign w2161 = w150 ~| w1740;
assign w2162 = w114 ~| w1741;
assign w2163 = w236 ~| w1741;
assign w2164 = w420 ~| w1742;
assign w2165 = w358 ~| w1742;
assign w2166 = w355 ~| w1743;
assign w2167 = w144 ~| w1743;
assign w2168 = w400 ~| w1744;
assign w2169 = w186 ~| w1744;
assign w2170 = w499 ~| w1745;
assign w2171 = w430 ~| w1745;
assign w2172 = w490 ~| w1746;
assign w2173 = w326 ~| w1746;
assign w2174 = w297 ~| w1747;
assign w2175 = w197 ~| w1747;
assign w2176 = w386 ~| w1748;
assign w2177 = w137 ~| w1748;
assign w2178 = w457 ~| w1749;
assign w2179 = w78 ~| w1749;
assign w2180 = w465 ~| w1750;
assign w2181 = w175 ~| w1750;
assign w2182 = w272 ~| w1751;
assign w2183 = w259 ~| w1751;
assign w2184 = w28 ~| w1752;
assign w2185 = w54 ~| w1752;
assign w2186 = w109 ~| w1753;
assign w2187 = w424 ~| w1754;
assign w2188 = w215 ~| w1754;
assign w2189 = w14 ~| w1755;
assign w2190 = w36 ~| w1755;
assign w2191 = w317 ~| w1756;
assign w2192 = w91 ~| w1756;
assign w2193 = w358 ~| w1757;
assign w2194 = w241 ~| w1757;
assign w2195 = w1470 | w1758;
assign w2196 = w70 ~| w1761;
assign w2197 = w90 ~| w1761;
assign w2198 = w124 ~| w1762;
assign w2199 = w196 ~| w1762;
assign w2200 = w457 ~| w1763;
assign w2201 = w414 ~| w1763;
assign w2202 = w106 ~| w1764;
assign w2203 = w214 ~| w1764;
assign w2204 = w268 ~| w1765;
assign w2205 = w240 ~| w1765;
assign w2206 = w487 ~| w1766;
assign w2207 = w381 ~| w1766;
assign w2208 = w29 ~| w1767;
assign w2209 = w264 ~| w1767;
assign w2210 = w472 ~| w1768;
assign w2211 = w1480 & w1768;
assign w2212 = w352 ~| w1769;
assign w2213 = w178 ~| w1769;
assign w2214 = w334 ~| w1770;
assign w2215 = w142 ~| w1770;
assign w2216 = w445 ~| w1771;
assign w2217 = w373 ~| w1771;
assign w2218 = w290 ~| w1772;
assign w2219 = w34 ~| w1772;
assign w2220 = w304 ~| w1773;
assign w2221 = w52 ~| w1773;
assign w2222 = w397 ~| w1774;
assign w2223 = w160 ~| w1774;
assign w2224 = w376 ~| w1775;
assign w2225 = w115 ~| w1775;
assign w2226 = w47 ~| w1776;
assign w2227 = w74 ~| w1776;
assign w2228 = w294 ~| w1777;
assign w2229 = w245 ~| w1777;
assign w2230 = w459 ~| w1778;
assign w2231 = w398 ~| w1778;
assign w2232 = w370 ~| w1779;
assign w2233 = w4 ~| w1779;
assign w2234 = w331 ~| w1780;
assign w2235 = w313 ~| w1780;
assign w2236 = w277 ~| w1781;
assign w2237 = w217 ~| w1781;
assign w2238 = w173 ~| w1782;
assign w2239 = w263 ~| w1783;
assign w2240 = w187 ~| w1783;
assign w2241 = w207 ~| w1784;
assign w2242 = w416 ~| w1785;
assign w2243 = w65 ~| w1785;
assign w2244 = w30 ~| w1786;
assign w2245 = w103 ~| w1786;
assign w2246 = w442 ~| w1787;
assign w2247 = w133 ~| w1787;
assign w2248 = w352 ~| w1788;
assign w2249 = w155 ~| w1788;
assign w2250 = w26 ~| w1789;
assign w2251 = w164 ~| w1789;
assign w2252 = w235 ~| w1790;
assign w2253 = w222 ~| w1790;
assign w2254 = w262 ~| w1791;
assign w2255 = w139 ~| w1791;
assign w2256 = w278 ~| w1792;
assign w2257 = w157 ~| w1793;
assign w2258 = w113 ~| w1793;
assign w2259 = w362 ~| w1794;
assign w2260 = w5 ~| w1794;
assign w2261 = w396 ~| w1795;
assign w2262 = w346 ~| w1795;
assign w2263 = w291 ~| w1796;
assign w2264 = w38 ~| w1796;
assign w2265 = w189 ~| w1797;
assign w2266 = w63 ~| w1797;
assign w2267 = w328 ~| w1798;
assign w2268 = w209 ~| w1798;
assign w2269 = w310 ~| w1799;
assign w2270 = w99 ~| w1799;
assign w2271 = w391 ~| w1800;
assign w2272 = w71 ~| w1800;
assign w2273 = w22 ~| w1804;
assign w2274 = w365 ~| w1804;
assign w2275 = w1527 & w1804;
assign w2276 = w48 ~| w1805;
assign w2277 = w84 ~| w1805;
assign w2278 = w426 ~| w1806;
assign w2279 = w280 ~| w1806;
assign w2280 = w437 ~| w1807;
assign w2281 = w118 ~| w1807;
assign w2282 = w244 ~| w1808;
assign w2283 = w66 ~| w1808;
assign w2284 = w228 ~| w1809;
assign w2285 = w156 ~| w1809;
assign w2286 = w316 ~| w1810;
assign w2287 = w210 ~| w1810;
assign w2288 = w326 ~| w1811;
assign w2289 = w138 ~| w1811;
assign w2290 = w406 ~| w1812;
assign w2291 = w344 ~| w1812;
assign w2292 = w102 ~| w1813;
assign w2293 = w192 ~| w1813;
assign w2294 = w296 ~| w1814;
assign w2295 = w174 ~| w1814;
assign w2296 = w384 ~| w1815;
assign w2297 = w255 ~| w1815;
assign w2298 = w308 ~| w1819;
assign w2299 = w184 ~| w1819;
assign w2300 = w94 ~| w1820;
assign w2301 = w110 ~| w1820;
assign w2302 = w17 ~| w1821;
assign w2303 = w130 ~| w1821;
assign w2304 = w350 ~| w1822;
assign w2305 = w273 ~| w1822;
assign w2306 = w379 ~| w1823;
assign w2307 = w220 ~| w1823;
assign w2308 = w238 ~| w1823;
assign w2309 = w288 ~| w1824;
assign w2310 = w258 ~| w1824;
assign w2311 = w202 ~| w1824;
assign w2312 = w76 ~| w1825;
assign w2313 = w166 ~| w1825;
assign w2314 = w368 ~| w1826;
assign w2315 = w332 ~| w1826;
assign w2316 = w40 ~| w1827;
assign w2317 = w148 ~| w1827;
assign w2318 = w58 ~| w1828;
assign w2319 = w1561 & w1828;
assign w2320 = w85 ~| w1829;
assign w2321 = w100 ~| w1829;
assign w2322 = w283 ~| w1830;
assign w2323 = w254 ~| w1830;
assign w2324 = w336 ~| w1831;
assign w2325 = w42 ~| w1831;
assign w2326 = w239 ~| w1832;
assign w2327 = w117 ~| w1832;
assign w2328 = w200 ~| w1833;
assign w2329 = w229 ~| w1833;
assign w2330 = w53 ~| w1833;
assign w2331 = w318 ~| w1834;
assign w2332 = w295 ~| w1834;
assign w2333 = w125 ~| w1834;
assign w2334 = w0 ~| w1835;
assign w2335 = w193 ~| w1835;
assign w2336 = w146 ~| w1835;
assign w2337 = w340 ~| w1836;
assign w2338 = w20 ~| w1836;
assign w2339 = w169 ~| w1836;
assign w2340 = w1848 | w1854;
assign w2341 = w1844 | w1855;
assign w2342 = w242 ~| w1857;
assign w2343 = w62 ~| w1857;
assign w2344 = w80 ~| w1858;
assign w2345 = w188 ~| w1858;
assign w2346 = w224 ~| w1859;
assign w2347 = w206 ~| w1859;
assign w2348 = w324 ~| w1860;
assign w2349 = w300 ~| w1860;
assign w2350 = w276 ~| w1861;
assign w2351 = w116 ~| w1861;
assign w2352 = w152 ~| w1861;
assign w2353 = w31 ~| w1862;
assign w2354 = w134 ~| w1862;
assign w2355 = w1570 & w1862;
assign w2356 = w170 ~| w1863;
assign w2357 = w314 ~| w1863;
assign w2358 = w44 ~| w1863;
assign w2359 = w252 ~| w1864;
assign w2360 = w98 ~| w1864;
assign w2361 = ~w1865;
assign w2362 = w1574 ~^ w1866;
assign w2363 = w542 ~| w1866;
assign w2364 = w542 & w1866;
assign w2365 = w1161 ~| w1867;
assign w2366 = w1132 & w1868;
assign w2367 = w825 ~| w1869;
assign w2368 = w1552 ~| w1869;
assign w2369 = w1285 ~| w1869;
assign w2370 = w1520 ~| w1869;
assign w2371 = w1488 ~| w1869;
assign w2372 = w1231 ~| w1869;
assign w2373 = w685 ~| w1869;
assign w2374 = w1443 ~| w1869;
assign w2375 = w1387 ~| w1869;
assign w2376 = w1568 ~| w1869;
assign w2377 = w1336 ~| w1869;
assign w2378 = w608 & w1870;
assign w2379 = in2[1] ~| w1871;
assign w2380 = in2[1] & w1871;
assign w2381 = w545 ~| w1872;
assign w2382 = w1873 ~^ in3[2];
assign w2383 = w1203 | w1875;
assign w2384 = w1211 | w1879;
assign w2385 = w3 | w1882;
assign w2386 = w1586 | w1894;
assign w2387 = w1584 | w1900;
assign w2388 = w1874 | w1905;
assign w2389 = w1208 | w1908;
assign w2390 = w1201 | w1909;
assign w2391 = w1206 | w1910;
assign w2392 = w1199 | w1911;
assign w2393 = w1223 | w1912;
assign w2394 = w1222 | w1913;
assign w2395 = w1204 | w1914;
assign w2396 = w1224 | w1916;
assign w2397 = w1213 | w1917;
assign w2398 = w1214 | w1918;
assign w2399 = w1229 | w1919;
assign w2400 = w1230 | w1920;
assign w2401 = w1225 | w1921;
assign w2402 = w1210 | w1922;
assign w2403 = w1219 | w1923;
assign w2404 = w1220 | w1924;
assign w2405 = w1221 | w1925;
assign w2406 = w1216 | w1926;
assign w2407 = w1215 | w1927;
assign w2408 = w1207 | w1928;
assign w2409 = w1209 | w1929;
assign w2410 = w1218 | w1930;
assign w2411 = w1876 | w1931;
assign w2412 = w1200 | w1932;
assign w2413 = w1226 | w1934;
assign w2414 = w1227 | w1935;
assign w2415 = w1228 | w1936;
assign w2416 = w1212 | w1937;
assign w2417 = w1202 | w1938;
assign w2418 = w1251 | w1940;
assign w2419 = w1255 | w1941;
assign w2420 = w1276 | w1942;
assign w2421 = w1254 | w1943;
assign w2422 = w1259 | w1944;
assign w2423 = w1261 | w1945;
assign w2424 = w1271 | w1946;
assign w2425 = w1281 | w1947;
assign w2426 = w1262 | w1948;
assign w2427 = w1270 | w1949;
assign w2428 = w1272 | w1950;
assign w2429 = w1257 | w1951;
assign w2430 = w1253 | w1952;
assign w2431 = w1256 | w1956;
assign w2432 = w1260 | w1957;
assign w2433 = w1279 | w1958;
assign w2434 = w1269 | w1959;
assign w2435 = w1273 | w1960;
assign w2436 = w1265 | w1962;
assign w2437 = w1277 | w1965;
assign w2438 = w1263 | w1966;
assign w2439 = w1266 | w1967;
assign w2440 = w1267 | w1968;
assign w2441 = w1275 | w1970;
assign w2442 = w1250 | w1972;
assign w2443 = w1258 | w1976;
assign w2444 = w0 | w1979;
assign w2445 = w1280 | w1982;
assign w2446 = w1264 | w1983;
assign w2447 = w1637 | w1987;
assign w2448 = w1252 | w1989;
assign w2449 = w1274 | w1994;
assign w2450 = w1971 ~| w1995;
assign w2451 = w1268 | w1998;
assign w2452 = w1635 | w2003;
assign w2453 = w1306 | w2005;
assign w2454 = w1332 | w2006;
assign w2455 = w1322 | w2007;
assign w2456 = w1313 | w2009;
assign w2457 = w1323 | w2010;
assign w2458 = w1304 | w2011;
assign w2459 = w1301 | w2012;
assign w2460 = w1308 | w2013;
assign w2461 = w1317 | w2014;
assign w2462 = w1311 | w2015;
assign w2463 = w1307 | w2016;
assign w2464 = w1324 | w2017;
assign w2465 = w1319 | w2019;
assign w2466 = w1310 | w2020;
assign w2467 = w1312 | w2021;
assign w2468 = w1321 | w2022;
assign w2469 = w1314 | w2023;
assign w2470 = w1302 | w2025;
assign w2471 = w1326 | w2029;
assign w2472 = w1318 | w2034;
assign w2473 = w1331 | w2035;
assign w2474 = w1305 | w2037;
assign w2475 = w1309 | w2041;
assign w2476 = w1303 | w2042;
assign w2477 = w13 | w2044;
assign w2478 = w1670 | w2046;
assign w2479 = w1327 | w2047;
assign w2480 = w1315 | w2048;
assign w2481 = w1330 | w2049;
assign w2482 = w1672 | w2050;
assign w2483 = w1329 | w2059;
assign w2484 = w2036 ~| w2060;
assign w2485 = w1316 | w2061;
assign w2486 = w1320 | w2062;
assign w2487 = w1328 | w2068;
assign w2488 = w1356 | w2069;
assign w2489 = w1359 | w2070;
assign w2490 = w1354 | w2071;
assign w2491 = w1353 | w2074;
assign w2492 = w1363 | w2075;
assign w2493 = w1364 | w2076;
assign w2494 = w1357 | w2077;
assign w2495 = w1378 | w2078;
assign w2496 = w1373 | w2082;
assign w2497 = w1379 | w2084;
assign w2498 = w1355 | w2086;
assign w2499 = w1375 | w2090;
assign w2500 = w1381 | w2092;
assign w2501 = w1365 | w2095;
assign w2502 = w1361 | w2096;
assign w2503 = w1369 | w2098;
assign w2504 = w2081 | w2102;
assign w2505 = w1705 | w2105;
assign w2506 = w1360 | w2106;
assign w2507 = w7 | w2109;
assign w2508 = w1377 | w2110;
assign w2509 = w1374 | w2114;
assign w2510 = w1382 | w2116;
assign w2511 = w1366 | w2117;
assign w2512 = w1380 | w2118;
assign w2513 = w1376 | w2120;
assign w2514 = w1383 | w2121;
assign w2515 = w1362 | w2122;
assign w2516 = w1707 | w2123;
assign w2517 = w2094 | w2126;
assign w2518 = w1371 | w2127;
assign w2519 = w2101 ~| w2130;
assign w2520 = w1358 | w2131;
assign w2521 = w1370 | w2132;
assign w2522 = w1368 | w2133;
assign w2523 = w1431 | w2135;
assign w2524 = w1420 | w2137;
assign w2525 = w5 | w2138;
assign w2526 = w1726 | w2141;
assign w2527 = w1414 | w2142;
assign w2528 = w1403 | w2143;
assign w2529 = w1724 | w2144;
assign w2530 = w1425 | w2146;
assign w2531 = w1421 | w2148;
assign w2532 = w1408 | w2149;
assign w2533 = w2134 ~| w2150;
assign w2534 = w1411 | w2152;
assign w2535 = w1410 | w2153;
assign w2536 = w1417 | w2154;
assign w2537 = w1432 | w2155;
assign w2538 = w1407 | w2156;
assign w2539 = w1405 | w2157;
assign w2540 = w1426 | w2158;
assign w2541 = w1427 | w2160;
assign w2542 = w1409 | w2164;
assign w2543 = w1418 | w2165;
assign w2544 = w1412 | w2166;
assign w2545 = w1406 | w2167;
assign w2546 = w2139 | w2172;
assign w2547 = w1404 | w2175;
assign w2548 = w1429 | w2177;
assign w2549 = w1415 | w2179;
assign w2550 = w1422 | w2181;
assign w2551 = w1416 | w2184;
assign w2552 = w1423 | w2185;
assign w2553 = w1430 | w2186;
assign w2554 = w1428 | w2190;
assign w2555 = w1424 | w2192;
assign w2556 = w1760 | w2196;
assign w2557 = w1458 | w2199;
assign w2558 = w1475 | w2200;
assign w2559 = w1465 | w2201;
assign w2560 = w1455 | w2203;
assign w2561 = w1453 | w2204;
assign w2562 = w1460 | w2205;
assign w2563 = w1463 | w2206;
assign w2564 = w1466 | w2207;
assign w2565 = w2195 ~| w2208;
assign w2566 = w1456 | w2209;
assign w2567 = w1451 | w2210;
assign w2568 = w15 | w2211;
assign w2569 = w1473 | w2212;
assign w2570 = w1450 | w2213;
assign w2571 = w1459 | w2215;
assign w2572 = w1457 | w2216;
assign w2573 = w1469 | w2217;
assign w2574 = w1454 | w2218;
assign w2575 = w1452 | w2219;
assign w2576 = w1461 | w2220;
assign w2577 = w1759 | w2221;
assign w2578 = w1464 | w2222;
assign w2579 = w1471 | w2223;
assign w2580 = w1468 | w2226;
assign w2581 = w1472 | w2227;
assign w2582 = w1467 | w2228;
assign w2583 = w1474 | w2243;
assign w2584 = w1476 | w2244;
assign w2585 = w1462 | w2245;
assign w2586 = w1801 | w2250;
assign w2587 = w1506 | w2252;
assign w2588 = w1494 | w2254;
assign w2589 = w1803 | w2264;
assign w2590 = w1497 | w2272;
assign w2591 = w1509 | w2273;
assign w2592 = w1505 | w2274;
assign w2593 = w8 | w2275;
assign w2594 = w1510 | w2276;
assign w2595 = w1514 | w2277;
assign w2596 = w1493 | w2278;
assign w2597 = w1511 | w2280;
assign w2598 = w1500 | w2282;
assign w2599 = w1502 | w2283;
assign w2600 = w1513 | w2284;
assign w2601 = w1504 | w2285;
assign w2602 = w1495 | w2286;
assign w2603 = w1508 | w2287;
assign w2604 = w1501 | w2288;
assign w2605 = w1516 | w2289;
assign w2606 = w1503 | w2290;
assign w2607 = w1512 | w2291;
assign w2608 = w1496 | w2292;
assign w2609 = w1498 | w2293;
assign w2610 = w1507 | w2295;
assign w2611 = w1499 | w2296;
assign w2612 = w1515 | w2297;
assign w2613 = w1532 | w2298;
assign w2614 = w1551 | w2299;
assign w2615 = w1544 | w2300;
assign w2616 = w1547 | w2301;
assign w2617 = w1531 | w2302;
assign w2618 = w1538 | w2303;
assign w2619 = w1542 | w2304;
assign w2620 = w1550 | w2305;
assign w2621 = w1548 | w2306;
assign w2622 = w1535 | w2309;
assign w2623 = w1540 | w2310;
assign w2624 = w1549 | w2311;
assign w2625 = w1546 | w2312;
assign w2626 = w1537 | w2313;
assign w2627 = w1534 | w2314;
assign w2628 = w1543 | w2315;
assign w2629 = w1533 | w2316;
assign w2630 = w1545 | w2317;
assign w2631 = w1536 | w2318;
assign w2632 = w11 | w2319;
assign w2633 = w1817 | w2325;
assign w2634 = w2308 | w2328;
assign w2635 = w1539 | w2335;
assign w2636 = w1816 | w2338;
assign w2637 = w1099 | w2342;
assign w2638 = w1092 | w2343;
assign w2639 = w1093 | w2344;
assign w2640 = w1088 | w2345;
assign w2641 = w1090 | w2346;
assign w2642 = w1084 | w2347;
assign w2643 = w1098 | w2348;
assign w2644 = w1091 | w2349;
assign w2645 = w1083 | w2350;
assign w2646 = w1086 | w2351;
assign w2647 = w1095 | w2352;
assign w2648 = w1094 | w2353;
assign w2649 = w1089 | w2354;
assign w2650 = w0 | w2355;
assign w2651 = w1837 | w2356;
assign w2652 = w1085 | w2357;
assign w2653 = w1082 | w2358;
assign w2654 = w1097 | w2359;
assign w2655 = w1096 | w2360;
assign w2656 = w1104 ~| w2364;
assign w2657 = w2365 ~^ in3[2];
assign w2658 = in3[2] ~| w2366;
assign w2659 = ~w2366;
assign w2660 = w1186 | w2367;
assign w2661 = w2330 | w2368;
assign w2662 = w1975 | w2369;
assign w2663 = w2266 | w2370;
assign w2664 = w2197 | w2371;
assign w2665 = w1885 | w2372;
assign w2666 = w1114 ~| w2373;
assign w2667 = w2136 | w2374;
assign w2668 = w2125 | w2375;
assign w2669 = w1853 | w2376;
assign w2670 = w2064 | w2377;
assign w2671 = w104 ~^ w2378;
assign w2672 = w105 | w2378;
assign w2673 = w544 ~| w2381;
assign w2674 = w2385 ~^ in3[5];
assign w2675 = w2388 ~^ in3[5];
assign w2676 = w2387 ~| w2394;
assign w2677 = w2386 ~| w2406;
assign w2678 = w2444 ~^ in3[8];
assign w2679 = w2429 ~| w2447;
assign w2680 = w2450 ~^ in3[8];
assign w2681 = w2419 ~| w2452;
assign w2682 = w2477 ~^ in3[11];
assign w2683 = w2454 ~| w2478;
assign w2684 = w2458 ~| w2482;
assign w2685 = w2484 ~^ in3[11];
assign w2686 = w2497 ~| w2505;
assign w2687 = w2507 ~^ in3[14];
assign w2688 = w2498 ~| w2516;
assign w2689 = w2519 ~^ in3[14];
assign w2690 = w2525 ~^ in3[17];
assign w2691 = w2533 ~^ in3[17];
assign w2692 = w2529 ~| w2551;
assign w2693 = w2526 ~| w2554;
assign w2694 = w2565 ~^ in3[20];
assign w2695 = w2568 ~^ in3[20];
assign w2696 = w2556 ~| w2580;
assign w2697 = w2577 ~| w2584;
assign w2698 = w1802 ~| w2591;
assign w2699 = w2593 ~^ in3[23];
assign w2700 = w2589 ~| w2595;
assign w2701 = w2586 ~| w2599;
assign w2702 = w1818 ~| w2617;
assign w2703 = w2632 ~^ in3[26];
assign w2704 = w2625 ~| w2633;
assign w2705 = w2631 ~| w2636;
assign w2706 = w2340 ~| w2638;
assign w2707 = w2341 ~| w2639;
assign w2708 = w1856 ~| w2648;
assign w2709 = w2650 ~^ in3[29];
assign w2710 = w2363 | w2656;
assign w2711 = ~w2657;
assign w2712 = w546 | w2659;
assign w2713 = w1140 ~| w2660;
assign w2714 = w2615 ~| w2661;
assign w2715 = w2418 ~| w2662;
assign w2716 = w2608 ~| w2663;
assign w2717 = w2583 ~| w2664;
assign w2718 = w2391 ~| w2665;
assign w2719 = w1130 & w2666;
assign w2720 = w2552 ~| w2667;
assign w2721 = w2493 ~| w2668;
assign w2722 = w2655 ~| w2669;
assign w2723 = w2469 ~| w2670;
assign w2724 = ~w2671;
assign w2725 = w1399 ~| w2671;
assign w2726 = w1245 ~| w2671;
assign w2727 = w1477 ~| w2671;
assign w2728 = w1295 ~| w2671;
assign w2729 = w1569 ~| w2671;
assign w2730 = w1348 ~| w2671;
assign w2731 = w1439 ~| w2671;
assign w2732 = w685 ~| w2671;
assign w2733 = w609 & w2672;
assign w2734 = w2379 ~| w2673;
assign w2735 = w549 ~^ w2674;
assign w2736 = w550 & w2674;
assign w2737 = w540 ~| w2675;
assign w2738 = ~w2675;
assign w2739 = w2676 ~^ in3[5];
assign w2740 = w2677 ~^ in3[5];
assign w2741 = w555 ~^ w2678;
assign w2742 = w556 & w2678;
assign w2743 = w2679 ~^ in3[8];
assign w2744 = w2680 ~^ in2[7];
assign w2745 = in2[7] & w2680;
assign w2746 = in2[7] | w2680;
assign w2747 = w2681 ~^ in3[8];
assign w2748 = w561 ~^ w2682;
assign w2749 = w562 & w2682;
assign w2750 = w2683 ~^ in3[11];
assign w2751 = w2684 ~^ in3[11];
assign w2752 = w2685 ~^ in2[10];
assign w2753 = in2[10] & w2685;
assign w2754 = in2[10] | w2685;
assign w2755 = w2686 ~^ in3[14];
assign w2756 = w567 ~^ w2687;
assign w2757 = w569 & w2687;
assign w2758 = w2688 ~^ in3[14];
assign w2759 = w2689 ~^ in2[13];
assign w2760 = in2[13] | w2689;
assign w2761 = in2[13] & w2689;
assign w2762 = w573 ~^ w2690;
assign w2763 = w574 & w2690;
assign w2764 = w2691 ~^ in2[16];
assign w2765 = in2[16] & w2691;
assign w2766 = in2[16] | w2691;
assign w2767 = w2692 ~^ in3[17];
assign w2768 = w2693 ~^ in3[17];
assign w2769 = w2694 ~^ in2[19];
assign w2770 = in2[19] & w2694;
assign w2771 = in2[19] | w2694;
assign w2772 = w579 ~^ w2695;
assign w2773 = w581 & w2695;
assign w2774 = w2696 ~^ in3[20];
assign w2775 = w2697 ~^ in3[20];
assign w2776 = w2698 ~^ in3[23];
assign w2777 = w585 ~^ w2699;
assign w2778 = w587 & w2699;
assign w2779 = w2700 ~^ in3[23];
assign w2780 = w2701 ~^ in3[23];
assign w2781 = w2702 ~^ in3[26];
assign w2782 = w591 ~^ w2703;
assign w2783 = w593 & w2703;
assign w2784 = w2704 ~^ in3[26];
assign w2785 = w2705 ~^ in3[26];
assign w2786 = w2706 ~^ in3[29];
assign w2787 = w2707 ~^ in3[29];
assign w2788 = w2708 ~^ in3[29];
assign w2789 = w597 ~^ w2709;
assign w2790 = w598 & w2709;
assign w2791 = ~w2712;
assign w2792 = w2713 ~^ in3[2];
assign w2793 = w2714 ~^ in3[26];
assign w2794 = w2715 ~^ in3[8];
assign w2795 = w2716 ~^ in3[23];
assign w2796 = w2717 ~^ in3[20];
assign w2797 = w2718 ~^ in3[5];
assign w2798 = ~w2719;
assign w2799 = w2720 ~^ in3[17];
assign w2800 = w2721 ~^ in3[14];
assign w2801 = w2722 ~^ in3[29];
assign w2802 = w2723 ~^ in3[11];
assign w2803 = ~w2724;
assign w2804 = w1068 & w2724;
assign w2805 = w2129 | w2725;
assign w2806 = w1886 | w2726;
assign w2807 = w2202 | w2727;
assign w2808 = w1991 | w2728;
assign w2809 = w1843 | w2729;
assign w2810 = w2052 | w2730;
assign w2811 = w2162 | w2731;
assign w2812 = w761 ~| w2732;
assign w2813 = w122 ~^ w2733;
assign w2814 = w123 | w2733;
assign w2815 = w2380 ~| w2734;
assign w2816 = w2382 & w2735;
assign w2817 = w2382 ~| w2735;
assign w2818 = w551 | w2736;
assign w2819 = in2[4] | w2738;
assign w2820 = w2739 ~^ w2741;
assign w2821 = w2739 | w2741;
assign w2822 = w2739 & w2741;
assign w2823 = w557 | w2742;
assign w2824 = w2747 ~^ w2748;
assign w2825 = w2747 | w2748;
assign w2826 = w2747 & w2748;
assign w2827 = w563 | w2749;
assign w2828 = w2750 ~^ w2756;
assign w2829 = w2750 | w2756;
assign w2830 = w2750 & w2756;
assign w2831 = w568 | w2757;
assign w2832 = w2755 ~^ w2762;
assign w2833 = w2755 & w2762;
assign w2834 = w2755 | w2762;
assign w2835 = w575 | w2763;
assign w2836 = w2767 ~^ w2772;
assign w2837 = w2767 | w2772;
assign w2838 = w2767 & w2772;
assign w2839 = w580 | w2773;
assign w2840 = w2776 ~^ in2[22];
assign w2841 = in2[22] | w2776;
assign w2842 = in2[22] & w2776;
assign w2843 = w2775 ~^ w2777;
assign w2844 = w2775 & w2777;
assign w2845 = w2775 | w2777;
assign w2846 = w586 | w2778;
assign w2847 = w2781 ~^ in2[25];
assign w2848 = in2[25] | w2781;
assign w2849 = in2[25] & w2781;
assign w2850 = w2780 ~^ w2782;
assign w2851 = w2780 | w2782;
assign w2852 = w2780 & w2782;
assign w2853 = w592 | w2783;
assign w2854 = w1103 ~^ w2786;
assign w2855 = w1103 | w2786;
assign w2856 = w1103 & w2786;
assign w2857 = w2362 ~^ w2787;
assign w2858 = w2362 & w2787;
assign w2859 = w2362 | w2787;
assign w2860 = w2788 ~^ in2[28];
assign w2861 = in2[28] | w2788;
assign w2862 = in2[28] & w2788;
assign w2863 = w2785 ~^ w2789;
assign w2864 = w2785 & w2789;
assign w2865 = w2785 | w2789;
assign w2866 = w599 | w2790;
assign w2867 = w2658 | w2791;
assign w2868 = ~w2791;
assign w2869 = ~w2798;
assign w2870 = w1560 ~| w2803;
assign w2871 = w837 ~| w2803;
assign w2872 = w2281 | w2804;
assign w2873 = w2489 ~| w2805;
assign w2874 = w2396 ~| w2806;
assign w2875 = w2581 ~| w2807;
assign w2876 = w2422 ~| w2808;
assign w2877 = w2646 ~| w2809;
assign w2878 = w2473 ~| w2810;
assign w2879 = w2549 ~| w2811;
assign w2880 = w1577 & w2812;
assign w2881 = w1489 ~| w2813;
assign w2882 = w1571 ~| w2813;
assign w2883 = w1343 ~| w2813;
assign w2884 = w1523 ~| w2813;
assign w2885 = w1394 ~| w2813;
assign w2886 = w1292 ~| w2813;
assign w2887 = w1558 ~| w2813;
assign w2888 = w1240 ~| w2813;
assign w2889 = w1441 ~| w2813;
assign w2890 = w832 ~| w2813;
assign w2891 = w685 ~| w2813;
assign w2892 = w610 & w2814;
assign w2893 = w2818 ~^ in2[4];
assign w2894 = w2818 & w2819;
assign w2895 = w2744 ~^ w2823;
assign w2896 = w2746 & w2823;
assign w2897 = w2752 ~^ w2827;
assign w2898 = w2754 & w2827;
assign w2899 = w2759 ~^ w2831;
assign w2900 = w2760 & w2831;
assign w2901 = w2764 ~^ w2835;
assign w2902 = w2766 & w2835;
assign w2903 = w2769 ~^ w2839;
assign w2904 = w2771 & w2839;
assign w2905 = w2840 ~^ w2846;
assign w2906 = w2841 & w2846;
assign w2907 = w2847 ~^ w2853;
assign w2908 = w2848 & w2853;
assign w2909 = w2860 ~^ w2866;
assign w2910 = w2861 & w2866;
assign w2911 = w2719 & w2868;
assign w2912 = w2712 ~^ w2869;
assign w2913 = w2712 | w2869;
assign w2914 = w2320 | w2870;
assign w2915 = w1188 | w2871;
assign w2916 = w2590 ~| w2872;
assign w2917 = w2873 ~^ in3[14];
assign w2918 = w2874 ~^ in3[5];
assign w2919 = w2875 ~^ in3[20];
assign w2920 = w2876 ~^ in3[8];
assign w2921 = w2877 ~^ in3[29];
assign w2922 = w2878 ~^ in3[11];
assign w2923 = w2879 ~^ in3[17];
assign w2924 = ~w2880;
assign w2925 = in3[5] & w2880;
assign w2926 = w2798 | w2880;
assign w2927 = w2198 | w2881;
assign w2928 = w1846 | w2882;
assign w2929 = w2054 | w2883;
assign w2930 = w2270 | w2884;
assign w2931 = w2103 | w2885;
assign w2932 = w1973 | w2886;
assign w2933 = w2321 | w2887;
assign w2934 = w1880 | w2888;
assign w2935 = w2147 | w2889;
assign w2936 = w1170 | w2890;
assign w2937 = w1111 ~| w2891;
assign w2938 = w140 ~^ w2892;
assign w2939 = w141 | w2892;
assign w2940 = w2675 ~^ w2893;
assign w2941 = w2737 | w2894;
assign w2942 = w2740 ~^ w2895;
assign w2943 = w2740 | w2895;
assign w2944 = w2740 & w2895;
assign w2945 = w2745 | w2896;
assign w2946 = w2743 ~^ w2897;
assign w2947 = w2743 | w2897;
assign w2948 = w2743 & w2897;
assign w2949 = w2753 | w2898;
assign w2950 = w2751 ~^ w2899;
assign w2951 = w2751 | w2899;
assign w2952 = w2751 & w2899;
assign w2953 = w2761 | w2900;
assign w2954 = w2758 ~^ w2901;
assign w2955 = w2758 & w2901;
assign w2956 = w2758 | w2901;
assign w2957 = w2765 | w2902;
assign w2958 = w2768 ~^ w2903;
assign w2959 = w2768 & w2903;
assign w2960 = w2768 | w2903;
assign w2961 = w2770 | w2904;
assign w2962 = w2774 ~^ w2905;
assign w2963 = w2774 | w2905;
assign w2964 = w2774 & w2905;
assign w2965 = w2842 | w2906;
assign w2966 = w2779 ~^ w2907;
assign w2967 = w2779 & w2907;
assign w2968 = w2779 | w2907;
assign w2969 = w2849 | w2908;
assign w2970 = w2784 ~^ w2909;
assign w2971 = w2784 | w2909;
assign w2972 = w2784 & w2909;
assign w2973 = w2862 | w2910;
assign w2974 = w2616 ~| w2914;
assign w2975 = w1148 ~| w2915;
assign w2976 = w2916 ~^ in3[23];
assign w2977 = w2719 ~| w2924;
assign w2978 = ~w2924;
assign w2979 = w2585 ~| w2927;
assign w2980 = w2649 ~| w2928;
assign w2981 = w2456 ~| w2929;
assign w2982 = w2605 ~| w2930;
assign w2983 = w2503 ~| w2931;
assign w2984 = w2433 ~| w2932;
assign w2985 = w2618 ~| w2933;
assign w2986 = w2395 ~| w2934;
assign w2987 = w2555 ~| w2935;
assign w2988 = w1136 ~| w2936;
assign w2989 = w1124 & w2937;
assign w2990 = w825 ~| w2938;
assign w2991 = w685 ~| w2938;
assign w2992 = w1336 ~| w2938;
assign w2993 = w1435 ~| w2938;
assign w2994 = w1387 ~| w2938;
assign w2995 = w1528 ~| w2938;
assign w2996 = w1558 ~| w2938;
assign w2997 = w1485 ~| w2938;
assign w2998 = w1231 ~| w2938;
assign w2999 = w1569 ~| w2938;
assign w3000 = w1285 ~| w2938;
assign w3001 = w611 & w2939;
assign w3002 = w2711 ~| w2940;
assign w3003 = ~w2940;
assign w3004 = w2974 ~^ in3[26];
assign w3005 = w2975 ~^ in3[2];
assign w3006 = w2719 ~^ w2978;
assign w3007 = in3[5] | w2978;
assign w3008 = w2979 ~^ in3[20];
assign w3009 = w2980 ~^ in3[29];
assign w3010 = w2981 ~^ in3[11];
assign w3011 = w2982 ~^ in3[23];
assign w3012 = w2983 ~^ in3[14];
assign w3013 = w2984 ~^ in3[8];
assign w3014 = w2985 ~^ in3[26];
assign w3015 = w2986 ~^ in3[5];
assign w3016 = w2987 ~^ in3[17];
assign w3017 = w2988 ~^ in3[2];
assign w3018 = w2989 ~^ in3[5];
assign w3019 = w2925 | w2989;
assign w3020 = w1172 | w2990;
assign w3021 = w1109 ~| w2991;
assign w3022 = w2038 | w2992;
assign w3023 = w2161 | w2993;
assign w3024 = w2112 | w2994;
assign w3025 = w2258 | w2995;
assign w3026 = w2327 | w2996;
assign w3027 = w2225 | w2997;
assign w3028 = w1892 | w2998;
assign w3029 = w1839 | w2999;
assign w3030 = w1993 | w3000;
assign w3031 = w158 ~^ w3001;
assign w3032 = w159 | w3001;
assign w3033 = w2657 ~| w3003;
assign w3034 = w2880 ~^ w3018;
assign w3035 = w3007 & w3019;
assign w3036 = w1144 ~| w3020;
assign w3037 = w1120 & w3021;
assign w3038 = w2464 ~| w3022;
assign w3039 = w2553 ~| w3023;
assign w3040 = w2495 ~| w3024;
assign w3041 = w2601 ~| w3025;
assign w3042 = w2630 ~| w3026;
assign w3043 = w2571 ~| w3027;
assign w3044 = w2417 ~| w3028;
assign w3045 = w2647 ~| w3029;
assign w3046 = w2438 ~| w3030;
assign w3047 = w1567 ~| w3031;
assign w3048 = w1490 ~| w3031;
assign w3049 = w1560 ~| w3031;
assign w3050 = w1443 ~| w3031;
assign w3051 = w1298 ~| w3031;
assign w3052 = w1246 ~| w3031;
assign w3053 = w838 ~| w3031;
assign w3054 = w1520 ~| w3031;
assign w3055 = w1400 ~| w3031;
assign w3056 = w685 ~| w3031;
assign w3057 = w1349 ~| w3031;
assign w3058 = w612 & w3032;
assign w3059 = ~w3034;
assign w3060 = ~w3035;
assign w3061 = w3036 ~^ in3[2];
assign w3062 = ~w3037;
assign w3063 = ~w3037;
assign w3064 = w3038 ~^ in3[11];
assign w3065 = w3039 ~^ in3[17];
assign w3066 = w3040 ~^ in3[14];
assign w3067 = w3041 ~^ in3[23];
assign w3068 = w3042 ~^ in3[26];
assign w3069 = w3043 ~^ in3[20];
assign w3070 = w3044 ~^ in3[5];
assign w3071 = w3045 ~^ in3[29];
assign w3072 = w3046 ~^ in3[8];
assign w3073 = w1087 | w3047;
assign w3074 = w2247 | w3048;
assign w3075 = w2333 | w3049;
assign w3076 = w2145 | w3050;
assign w3077 = w1977 | w3051;
assign w3078 = w1878 | w3052;
assign w3079 = w1180 | w3053;
assign w3080 = w2255 | w3054;
assign w3081 = w2113 | w3055;
assign w3082 = w1119 ~| w3056;
assign w3083 = w2056 | w3057;
assign w3084 = w176 ~^ w3058;
assign w3085 = w177 | w3058;
assign w3086 = w3035 ~| w3062;
assign w3087 = ~w3063;
assign w3088 = w3035 ^ w3063;
assign w3089 = w2912 ~^ w3071;
assign w3090 = w2913 & w3071;
assign w3091 = w2651 ~| w3073;
assign w3092 = w2579 ~| w3074;
assign w3093 = w2626 ~| w3075;
assign w3094 = w2548 ~| w3076;
assign w3095 = w2426 ~| w3077;
assign w3096 = w2412 ~| w3078;
assign w3097 = w1138 ~| w3079;
assign w3098 = w2610 ~| w3080;
assign w3099 = w2502 ~| w3081;
assign w3100 = w1129 & w3082;
assign w3101 = w2460 ~| w3083;
assign w3102 = w1487 ~| w3084;
assign w3103 = w1555 ~| w3084;
assign w3104 = w831 ~| w3084;
assign w3105 = w1521 ~| w3084;
assign w3106 = w1393 ~| w3084;
assign w3107 = w1436 ~| w3084;
assign w3108 = w685 ~| w3084;
assign w3109 = w1291 ~| w3084;
assign w3110 = w1239 ~| w3084;
assign w3111 = w1572 ~| w3084;
assign w3112 = w1342 ~| w3084;
assign w3113 = w613 & w3085;
assign w3114 = w3060 | w3087;
assign w3115 = w2911 | w3090;
assign w3116 = w3091 ~^ in3[29];
assign w3117 = w3092 ~^ in3[20];
assign w3118 = w3093 ~^ in3[26];
assign w3119 = w3094 ~^ in3[17];
assign w3120 = w3095 ~^ in3[8];
assign w3121 = w3096 ~^ in3[5];
assign w3122 = w3097 ~^ in3[2];
assign w3123 = w3098 ~^ in3[23];
assign w3124 = w3099 ~^ in3[14];
assign w3125 = ~w3100;
assign w3126 = in3[8] | w3100;
assign w3127 = w3062 | w3100;
assign w3128 = w3101 ~^ in3[11];
assign w3129 = w2249 | w3102;
assign w3130 = w2336 | w3103;
assign w3131 = w1198 | w3104;
assign w3132 = w2257 | w3105;
assign w3133 = w2111 | w3106;
assign w3134 = w2140 | w3107;
assign w3135 = w1118 ~| w3108;
assign w3136 = w1981 | w3109;
assign w3137 = w1888 | w3110;
assign w3138 = w1849 | w3111;
assign w3139 = w2058 | w3112;
assign w3140 = w194 ~^ w3113;
assign w3141 = w195 | w3113;
assign w3142 = ~w3115;
assign w3143 = w3006 ~^ w3116;
assign w3144 = w2926 & w3116;
assign w3145 = w3037 ~| w3125;
assign w3146 = ~w3125;
assign w3147 = w2570 ~| w3129;
assign w3148 = w2614 ~| w3130;
assign w3149 = w1160 ~| w3131;
assign w3150 = w2609 ~| w3132;
assign w3151 = w2501 ~| w3133;
assign w3152 = w2545 ~| w3134;
assign w3153 = w1127 & w3135;
assign w3154 = w2440 ~| w3136;
assign w3155 = w2416 ~| w3137;
assign w3156 = w2640 ~| w3138;
assign w3157 = w2471 ~| w3139;
assign w3158 = w1441 ~| w3140;
assign w3159 = w1232 ~| w3140;
assign w3160 = w1286 ~| w3140;
assign w3161 = w1559 ~| w3140;
assign w3162 = w1337 ~| w3140;
assign w3163 = w826 ~| w3140;
assign w3164 = w685 ~| w3140;
assign w3165 = w1526 ~| w3140;
assign w3166 = w1487 ~| w3140;
assign w3167 = w1572 ~| w3140;
assign w3168 = w1388 ~| w3140;
assign w3169 = w614 & w3141;
assign w3170 = w3115 ~^ w3143;
assign w3171 = w3142 ~| w3143;
assign w3172 = ~w3143;
assign w3173 = w2977 | w3144;
assign w3174 = w3087 ~^ w3146;
assign w3175 = in3[8] & w3146;
assign w3176 = w3147 ~^ in3[20];
assign w3177 = w3148 ~^ in3[26];
assign w3178 = w3149 ~^ in3[2];
assign w3179 = w3150 ~^ in3[23];
assign w3180 = w3151 ~^ in3[14];
assign w3181 = w3152 ~^ in3[17];
assign w3182 = w3153 ~^ in3[8];
assign w3183 = w3154 ~^ in3[8];
assign w3184 = w3155 ~^ in3[5];
assign w3185 = w3156 ~^ in3[29];
assign w3186 = w3157 ~^ in3[11];
assign w3187 = w2151 | w3158;
assign w3188 = w1906 | w3159;
assign w3189 = w1985 | w3160;
assign w3190 = w2339 | w3161;
assign w3191 = w2040 | w3162;
assign w3192 = w1168 | w3163;
assign w3193 = w1115 ~| w3164;
assign w3194 = w2251 | w3165;
assign w3195 = w2238 | w3166;
assign w3196 = w1847 | w3167;
assign w3197 = w2115 | w3168;
assign w3198 = w212 ~^ w3169;
assign w3199 = w213 | w3169;
assign w3200 = w3115 | w3172;
assign w3201 = w3153 | w3175;
assign w3202 = w3100 ~^ w3182;
assign w3203 = w3034 ~^ w3185;
assign w3204 = w3059 | w3185;
assign w3205 = ~w3185;
assign w3206 = w2550 ~| w3187;
assign w3207 = w2399 ~| w3188;
assign w3208 = w2435 ~| w3189;
assign w3209 = w2624 ~| w3190;
assign w3210 = w2472 ~| w3191;
assign w3211 = w1156 ~| w3192;
assign w3212 = w1122 & w3193;
assign w3213 = w2603 ~| w3194;
assign w3214 = w2557 ~| w3195;
assign w3215 = w2642 ~| w3196;
assign w3216 = w2499 ~| w3197;
assign w3217 = w1440 ~| w3198;
assign w3218 = w1244 ~| w3198;
assign w3219 = w1478 ~| w3198;
assign w3220 = w1565 ~| w3198;
assign w3221 = w1555 ~| w3198;
assign w3222 = w1524 ~| w3198;
assign w3223 = w685 ~| w3198;
assign w3224 = w1347 ~| w3198;
assign w3225 = w836 ~| w3198;
assign w3226 = w1294 ~| w3198;
assign w3227 = w1398 ~| w3198;
assign w3228 = w615 & w3199;
assign w3229 = w3126 & w3201;
assign w3230 = ~w3202;
assign w3231 = w3173 ~^ w3203;
assign w3232 = w3173 & w3204;
assign w3233 = w3034 ~| w3205;
assign w3234 = w3206 ~^ in3[17];
assign w3235 = w3207 ~^ in3[5];
assign w3236 = w3208 ~^ in3[8];
assign w3237 = w3209 ~^ in3[26];
assign w3238 = w3210 ~^ in3[11];
assign w3239 = w3211 ~^ in3[2];
assign w3240 = ~w3212;
assign w3241 = ~w3212;
assign w3242 = w3213 ~^ in3[23];
assign w3243 = w3214 ~^ in3[20];
assign w3244 = w3215 ~^ in3[29];
assign w3245 = w3216 ~^ in3[14];
assign w3246 = w2169 | w3217;
assign w3247 = w1896 | w3218;
assign w3248 = w2240 | w3219;
assign w3249 = w1842 | w3220;
assign w3250 = w2307 | w3221;
assign w3251 = w2265 | w3222;
assign w3252 = w1107 ~| w3223;
assign w3253 = w2066 | w3224;
assign w3254 = w1177 | w3225;
assign w3255 = w1986 | w3226;
assign w3256 = w2119 | w3227;
assign w3257 = w230 ~^ w3228;
assign w3258 = w231 | w3228;
assign w3259 = ~w3229;
assign w3260 = ~w3231;
assign w3261 = w3232 | w3233;
assign w3262 = w3229 ~| w3240;
assign w3263 = ~w3241;
assign w3264 = w3229 ^ w3241;
assign w3265 = w3088 ~^ w3244;
assign w3266 = w3114 & w3244;
assign w3267 = w2532 ~| w3246;
assign w3268 = w2389 ~| w3247;
assign w3269 = w2560 ~| w3248;
assign w3270 = w2641 ~| w3249;
assign w3271 = w2635 ~| w3250;
assign w3272 = w2600 ~| w3251;
assign w3273 = w1128 & w3252;
assign w3274 = w2466 ~| w3253;
assign w3275 = w1154 ~| w3254;
assign w3276 = w2420 ~| w3255;
assign w3277 = w2491 ~| w3256;
assign w3278 = w828 ~| w3257;
assign w3279 = w1557 ~| w3257;
assign w3280 = w1288 ~| w3257;
assign w3281 = w1236 ~| w3257;
assign w3282 = w1339 ~| w3257;
assign w3283 = w1438 ~| w3257;
assign w3284 = w685 ~| w3257;
assign w3285 = w1390 ~| w3257;
assign w3286 = w1525 ~| w3257;
assign w3287 = w1571 ~| w3257;
assign w3288 = w1479 ~| w3257;
assign w3289 = w616 & w3258;
assign w3290 = ~w3261;
assign w3291 = w3259 | w3263;
assign w3292 = w3261 ~^ w3265;
assign w3293 = ~w3265;
assign w3294 = w3086 | w3266;
assign w3295 = w3267 ~^ in3[17];
assign w3296 = w3268 ~^ in3[5];
assign w3297 = w3269 ~^ in3[20];
assign w3298 = w3270 ~^ in3[29];
assign w3299 = w3271 ~^ in3[26];
assign w3300 = w3272 ~^ in3[23];
assign w3301 = ~w3273;
assign w3302 = in3[11] | w3273;
assign w3303 = w3240 | w3273;
assign w3304 = w3274 ~^ in3[11];
assign w3305 = w3275 ~^ in3[2];
assign w3306 = w3276 ~^ in3[8];
assign w3307 = w3277 ~^ in3[14];
assign w3308 = w1176 | w3278;
assign w3309 = w1541 | w3279;
assign w3310 = w1997 | w3280;
assign w3311 = w1884 | w3281;
assign w3312 = w2051 | w3282;
assign w3313 = w2163 | w3283;
assign w3314 = w1117 ~| w3284;
assign w3315 = w2107 | w3285;
assign w3316 = w2268 | w3286;
assign w3317 = w1840 | w3287;
assign w3318 = w2241 | w3288;
assign w3319 = w248 ~^ w3289;
assign w3320 = w249 | w3289;
assign w3321 = w3265 ~| w3290;
assign w3322 = w3261 | w3293;
assign w3323 = ~w3294;
assign w3324 = w3174 ~^ w3298;
assign w3325 = w3127 & w3298;
assign w3326 = w3170 ~^ w3299;
assign w3327 = w3200 & w3299;
assign w3328 = w3212 ~| w3301;
assign w3329 = ~w3301;
assign w3330 = w1142 ~| w3308;
assign w3331 = w2634 ~| w3309;
assign w3332 = w2430 ~| w3310;
assign w3333 = w2400 ~| w3311;
assign w3334 = w2470 ~| w3312;
assign w3335 = w2547 ~| w3313;
assign w3336 = w1121 & w3314;
assign w3337 = w2494 ~| w3315;
assign w3338 = w2598 ~| w3316;
assign w3339 = w2637 ~| w3317;
assign w3340 = w2562 ~| w3318;
assign w3341 = w1235 ~| w3319;
assign w3342 = w1338 ~| w3319;
assign w3343 = w685 ~| w3319;
assign w3344 = w827 ~| w3319;
assign w3345 = w1389 ~| w3319;
assign w3346 = w1437 ~| w3319;
assign w3347 = w1553 ~| w3319;
assign w3348 = w1479 ~| w3319;
assign w3349 = w1527 ~| w3319;
assign w3350 = w1570 ~| w3319;
assign w3351 = w1287 ~| w3319;
assign w3352 = w617 & w3320;
assign w3353 = w3294 ~^ w3324;
assign w3354 = w3323 ~| w3324;
assign w3355 = ~w3324;
assign w3356 = w3145 | w3325;
assign w3357 = ~w3326;
assign w3358 = w3171 | w3327;
assign w3359 = w3263 ~^ w3329;
assign w3360 = in3[11] & w3329;
assign w3361 = w3330 ~^ in3[2];
assign w3362 = w3331 ~^ in3[26];
assign w3363 = w3332 ~^ in3[8];
assign w3364 = w3333 ~^ in3[5];
assign w3365 = w3334 ~^ in3[11];
assign w3366 = w3335 ~^ in3[17];
assign w3367 = w3336 ~^ in3[11];
assign w3368 = w3337 ~^ in3[14];
assign w3369 = w3338 ~^ in3[23];
assign w3370 = w3339 ~^ in3[29];
assign w3371 = w3340 ~^ in3[20];
assign w3372 = w1881 | w3341;
assign w3373 = w2043 | w3342;
assign w3374 = w1112 ~| w3343;
assign w3375 = w1173 | w3344;
assign w3376 = w2108 | w3345;
assign w3377 = w2188 | w3346;
assign w3378 = w2329 | w3347;
assign w3379 = w2237 | w3348;
assign w3380 = w2253 | w3349;
assign w3381 = w1845 | w3350;
assign w3382 = w1978 | w3351;
assign w3383 = w266 ~^ w3352;
assign w3384 = w267 | w3352;
assign w3385 = w3294 | w3355;
assign w3386 = w3336 | w3360;
assign w3387 = w3231 ~^ w3362;
assign w3388 = w3260 | w3362;
assign w3389 = ~w3362;
assign w3390 = w3273 ~^ w3367;
assign w3391 = w3202 ~^ w3370;
assign w3392 = w3230 | w3370;
assign w3393 = ~w3370;
assign w3394 = w2393 ~| w3372;
assign w3395 = w2453 ~| w3373;
assign w3396 = w1126 & w3374;
assign w3397 = w1163 ~| w3375;
assign w3398 = w2500 ~| w3376;
assign w3399 = w2531 ~| w3377;
assign w3400 = w2623 ~| w3378;
assign w3401 = w2566 ~| w3379;
assign w3402 = w2612 ~| w3380;
assign w3403 = w2654 ~| w3381;
assign w3404 = w2437 ~| w3382;
assign w3405 = w1391 ~| w3383;
assign w3406 = w1445 ~| w3383;
assign w3407 = w1519 ~| w3383;
assign w3408 = w1569 ~| w3383;
assign w3409 = w829 ~| w3383;
assign w3410 = w1289 ~| w3383;
assign w3411 = w1486 ~| w3383;
assign w3412 = w685 ~| w3383;
assign w3413 = w1552 ~| w3383;
assign w3414 = w1340 ~| w3383;
assign w3415 = w1237 ~| w3383;
assign w3416 = w618 & w3384;
assign w3417 = w3302 & w3386;
assign w3418 = w3358 ~^ w3387;
assign w3419 = w3358 & w3388;
assign w3420 = w3231 ~| w3389;
assign w3421 = ~w3390;
assign w3422 = w3356 ~^ w3391;
assign w3423 = w3356 & w3392;
assign w3424 = w3202 ~| w3393;
assign w3425 = w3394 ~^ in3[5];
assign w3426 = w3395 ~^ in3[11];
assign w3427 = ~w3396;
assign w3428 = w3397 ~^ in3[2];
assign w3429 = w3398 ~^ in3[14];
assign w3430 = w3399 ~^ in3[17];
assign w3431 = w3400 ~^ in3[26];
assign w3432 = w3401 ~^ in3[20];
assign w3433 = w3402 ~^ in3[23];
assign w3434 = w3403 ~^ in3[29];
assign w3435 = w3404 ~^ in3[8];
assign w3436 = w2104 | w3405;
assign w3437 = w2194 | w3406;
assign w3438 = w2279 | w3407;
assign w3439 = w1841 | w3408;
assign w3440 = w1197 | w3409;
assign w3441 = w1988 | w3410;
assign w3442 = w2229 | w3411;
assign w3443 = w1116 | w3412;
assign w3444 = w2326 | w3413;
assign w3445 = w2057 | w3414;
assign w3446 = w1877 | w3415;
assign w3447 = w284 ~^ w3416;
assign w3448 = w285 | w3416;
assign w3449 = w3396 ~^ w3417;
assign w3450 = ~w3417;
assign w3451 = ~w3418;
assign w3452 = w3419 | w3420;
assign w3453 = ~w3422;
assign w3454 = w3423 | w3424;
assign w3455 = w3417 ~| w3427;
assign w3456 = ~w3427;
assign w3457 = w3292 ~^ w3431;
assign w3458 = w3322 & w3431;
assign w3459 = w3264 ~^ w3434;
assign w3460 = w3291 & w3434;
assign w3461 = w2496 ~| w3436;
assign w3462 = w2524 ~| w3437;
assign w3463 = w2587 ~| w3438;
assign w3464 = w2645 ~| w3439;
assign w3465 = w1153 ~| w3440;
assign w3466 = w2424 ~| w3441;
assign w3467 = w2561 ~| w3442;
assign w3468 = w1125 ~| w3443;
assign w3469 = w2620 ~| w3444;
assign w3470 = w2455 ~| w3445;
assign w3471 = w2408 ~| w3446;
assign w3472 = w1567 ~| w3447;
assign w3473 = w1522 ~| w3447;
assign w3474 = w823 ~| w3447;
assign w3475 = w1334 ~| w3447;
assign w3476 = w1385 ~| w3447;
assign w3477 = w1481 ~| w3447;
assign w3478 = w1233 ~| w3447;
assign w3479 = w1283 ~| w3447;
assign w3480 = w1557 ~| w3447;
assign w3481 = w1444 ~| w3447;
assign w3482 = w619 & w3448;
assign w3483 = ~w3452;
assign w3484 = ~w3454;
assign w3485 = w3450 | w3456;
assign w3486 = w3452 ~^ w3457;
assign w3487 = ~w3457;
assign w3488 = w3321 | w3458;
assign w3489 = w3454 ~^ w3459;
assign w3490 = ~w3459;
assign w3491 = w3262 | w3460;
assign w3492 = w3461 ~^ in3[14];
assign w3493 = w3462 ~^ in3[17];
assign w3494 = w3463 ~^ in3[23];
assign w3495 = w3464 ~^ in3[29];
assign w3496 = w3465 ~^ in3[2];
assign w3497 = w3466 ~^ in3[8];
assign w3498 = w3467 ~^ in3[20];
assign w3499 = w3456 ~^ w3468;
assign w3500 = w3469 ~^ in3[26];
assign w3501 = w3470 ~^ in3[11];
assign w3502 = w3471 ~^ in3[5];
assign w3503 = w1838 | w3472;
assign w3504 = w2294 | w3473;
assign w3505 = w1185 | w3474;
assign w3506 = w2039 | w3475;
assign w3507 = w2128 | w3476;
assign w3508 = w2239 | w3477;
assign w3509 = w1893 | w3478;
assign w3510 = w1974 | w3479;
assign w3511 = w2323 | w3480;
assign w3512 = w2183 | w3481;
assign w3513 = w302 ~^ w3482;
assign w3514 = w303 | w3482;
assign w3515 = w3457 ~| w3483;
assign w3516 = w3459 ~| w3484;
assign w3517 = w3452 | w3487;
assign w3518 = ~w3488;
assign w3519 = w3454 | w3490;
assign w3520 = ~w3491;
assign w3521 = w3359 ~^ w3495;
assign w3522 = w3303 & w3495;
assign w3523 = w3353 ~^ w3500;
assign w3524 = w3385 & w3500;
assign w3525 = w2644 ~| w3503;
assign w3526 = w2588 ~| w3504;
assign w3527 = w1147 ~| w3505;
assign w3528 = w2463 ~| w3506;
assign w3529 = w2490 ~| w3507;
assign w3530 = w2574 ~| w3508;
assign w3531 = w2404 ~| w3509;
assign w3532 = w2431 ~| w3510;
assign w3533 = w2622 ~| w3511;
assign w3534 = w2539 ~| w3512;
assign w3535 = w1335 ~| w3513;
assign w3536 = w1565 ~| w3513;
assign w3537 = w1529 ~| w3513;
assign w3538 = w1234 ~| w3513;
assign w3539 = w824 ~| w3513;
assign w3540 = w1284 ~| w3513;
assign w3541 = w1554 ~| w3513;
assign w3542 = w1482 ~| w3513;
assign w3543 = w1386 ~| w3513;
assign w3544 = w1446 ~| w3513;
assign w3545 = w620 & w3514;
assign w3546 = w3491 ~^ w3521;
assign w3547 = w3520 ~| w3521;
assign w3548 = ~w3521;
assign w3549 = w3328 | w3522;
assign w3550 = w3488 ~^ w3523;
assign w3551 = w3518 ~| w3523;
assign w3552 = ~w3523;
assign w3553 = w3354 | w3524;
assign w3554 = w3525 ~^ in3[29];
assign w3555 = w3526 ~^ in3[23];
assign w3556 = w3527 ~^ in3[2];
assign w3557 = w3528 ~^ in3[11];
assign w3558 = w3529 ~^ in3[14];
assign w3559 = w3530 ~^ in3[20];
assign w3560 = w3531 ~^ in3[5];
assign w3561 = w3532 ~^ in3[8];
assign w3562 = w3533 ~^ in3[26];
assign w3563 = w3534 ~^ in3[17];
assign w3564 = w2063 | w3535;
assign w3565 = w1851 | w3536;
assign w3566 = w2256 | w3537;
assign w3567 = w1887 | w3538;
assign w3568 = w1179 | w3539;
assign w3569 = w2002 | w3540;
assign w3570 = w2322 | w3541;
assign w3571 = w2236 | w3542;
assign w3572 = w2124 | w3543;
assign w3573 = w2182 | w3544;
assign w3574 = w320 ~^ w3545;
assign w3575 = w321 | w3545;
assign w3576 = w3491 | w3548;
assign w3577 = w3488 | w3552;
assign w3578 = w3390 ~^ w3554;
assign w3579 = w3421 | w3554;
assign w3580 = ~w3554;
assign w3581 = w3418 ~^ w3555;
assign w3582 = w3451 | w3555;
assign w3583 = ~w3555;
assign w3584 = w3422 ~^ w3562;
assign w3585 = w3453 | w3562;
assign w3586 = ~w3562;
assign w3587 = w2467 ~| w3564;
assign w3588 = w2652 ~| w3565;
assign w3589 = w2602 ~| w3566;
assign w3590 = w2390 ~| w3567;
assign w3591 = w1137 ~| w3568;
assign w3592 = w2423 ~| w3569;
assign w3593 = w2613 ~| w3570;
assign w3594 = w2576 ~| w3571;
assign w3595 = w2492 ~| w3572;
assign w3596 = w2541 ~| w3573;
assign w3597 = w1478 ~| w3574;
assign w3598 = w1568 ~| w3574;
assign w3599 = w1529 ~| w3574;
assign w3600 = w1296 ~| w3574;
assign w3601 = w1345 ~| w3574;
assign w3602 = w1242 ~| w3574;
assign w3603 = w1556 ~| w3574;
assign w3604 = w1396 ~| w3574;
assign w3605 = w1434 ~| w3574;
assign w3606 = w834 ~| w3574;
assign w3607 = w621 & w3575;
assign w3608 = w3549 ~^ w3578;
assign w3609 = w3549 & w3579;
assign w3610 = w3390 ~| w3580;
assign w3611 = w3418 ~| w3583;
assign w3612 = w3553 ~^ w3584;
assign w3613 = w3553 & w3585;
assign w3614 = w3422 ~| w3586;
assign w3615 = w3587 ~^ in3[11];
assign w3616 = w3588 ~^ in3[29];
assign w3617 = w3589 ~^ in3[23];
assign w3618 = w3590 ~^ in3[5];
assign w3619 = w3591 ~^ in3[2];
assign w3620 = w3592 ~^ in3[8];
assign w3621 = w3593 ~^ in3[26];
assign w3622 = w3594 ~^ in3[20];
assign w3623 = w3595 ~^ in3[14];
assign w3624 = w3596 ~^ in3[17];
assign w3625 = w2214 | w3597;
assign w3626 = w1850 | w3598;
assign w3627 = w2263 | w3599;
assign w3628 = w1990 | w3600;
assign w3629 = w2055 | w3601;
assign w3630 = w1899 | w3602;
assign w3631 = w2332 | w3603;
assign w3632 = w2091 | w3604;
assign w3633 = w2174 | w3605;
assign w3634 = w1191 | w3606;
assign w3635 = w338 ~^ w3607;
assign w3636 = w339 | w3607;
assign w3637 = ~w3608;
assign w3638 = w3609 | w3610;
assign w3639 = ~w3612;
assign w3640 = w3613 | w3614;
assign w3641 = w3449 ~^ w3616;
assign w3642 = w3485 & w3616;
assign w3643 = w3486 ~^ w3617;
assign w3644 = w3517 & w3617;
assign w3645 = w3489 ~^ w3621;
assign w3646 = w3519 & w3621;
assign w3647 = w2582 ~| w3625;
assign w3648 = w2643 ~| w3626;
assign w3649 = w2604 ~| w3627;
assign w3650 = w2428 ~| w3628;
assign w3651 = w2457 ~| w3629;
assign w3652 = w2398 ~| w3630;
assign w3653 = w2628 ~| w3631;
assign w3654 = w2509 ~| w3632;
assign w3655 = w2538 ~| w3633;
assign w3656 = w1146 ~| w3634;
assign w3657 = w1238 ~| w3635;
assign w3658 = w830 ~| w3635;
assign w3659 = w1392 ~| w3635;
assign w3660 = w1442 ~| w3635;
assign w3661 = w1290 ~| w3635;
assign w3662 = w1553 ~| w3635;
assign w3663 = w1341 ~| w3635;
assign w3664 = w1477 ~| w3635;
assign w3665 = w1523 ~| w3635;
assign w3666 = w622 & w3636;
assign w3667 = ~w3638;
assign w3668 = ~w3640;
assign w3669 = w3638 ~^ w3641;
assign w3670 = ~w3641;
assign w3671 = w3455 | w3642;
assign w3672 = ~w3643;
assign w3673 = w3515 | w3644;
assign w3674 = w3640 ~^ w3645;
assign w3675 = ~w3645;
assign w3676 = w3516 | w3646;
assign w3677 = w3647 ~^ in3[20];
assign w3678 = w3648 ~^ in3[29];
assign w3679 = w3649 ~^ in3[23];
assign w3680 = w3650 ~^ in3[8];
assign w3681 = w3651 ~^ in3[11];
assign w3682 = w3652 ~^ in3[5];
assign w3683 = w3653 ~^ in3[26];
assign w3684 = w3654 ~^ in3[14];
assign w3685 = w3655 ~^ in3[17];
assign w3686 = w3656 ~^ in3[2];
assign w3687 = w1891 | w3657;
assign w3688 = w1183 | w3658;
assign w3689 = w2083 | w3659;
assign w3690 = w2191 | w3660;
assign w3691 = w1980 | w3661;
assign w3692 = w2331 | w3662;
assign w3693 = w2045 | w3663;
assign w3694 = w2235 | w3664;
assign w3695 = w2269 | w3665;
assign w3696 = w356 ~^ w3666;
assign w3697 = w357 | w3666;
assign w3698 = w3641 ~| w3667;
assign w3699 = w3645 ~| w3668;
assign w3700 = w3638 | w3670;
assign w3701 = ~w3673;
assign w3702 = w3640 | w3675;
assign w3703 = ~w3676;
assign w3704 = w3499 ~^ w3678;
assign w3705 = w3550 ~^ w3679;
assign w3706 = w3577 & w3679;
assign w3707 = w3546 ~^ w3683;
assign w3708 = w3576 & w3683;
assign w3709 = w2405 ~| w3687;
assign w3710 = w1162 ~| w3688;
assign w3711 = w2515 ~| w3689;
assign w3712 = w2527 ~| w3690;
assign w3713 = w2432 ~| w3691;
assign w3714 = w2619 ~| w3692;
assign w3715 = w2462 ~| w3693;
assign w3716 = w2569 ~| w3694;
assign w3717 = w2607 ~| w3695;
assign w3718 = w1341 ~| w3696;
assign w3719 = w1518 ~| w3696;
assign w3720 = w1392 ~| w3696;
assign w3721 = w1435 ~| w3696;
assign w3722 = w1290 ~| w3696;
assign w3723 = w1561 ~| w3696;
assign w3724 = w1481 ~| w3696;
assign w3725 = w830 ~| w3696;
assign w3726 = w1238 ~| w3696;
assign w3727 = w623 & w3697;
assign w3728 = w3671 ~^ w3704;
assign w3729 = w3673 ~^ w3705;
assign w3730 = w3701 ~| w3705;
assign w3731 = ~w3705;
assign w3732 = w3551 | w3706;
assign w3733 = w3676 ~^ w3707;
assign w3734 = w3703 ~| w3707;
assign w3735 = ~w3707;
assign w3736 = w3547 | w3708;
assign w3737 = w3709 ~^ in3[5];
assign w3738 = w3710 ~^ in3[2];
assign w3739 = w3711 ~^ in3[14];
assign w3740 = w3712 ~^ in3[17];
assign w3741 = w3713 ~^ in3[8];
assign w3742 = w3714 ~^ in3[26];
assign w3743 = w3715 ~^ in3[11];
assign w3744 = w3716 ~^ in3[20];
assign w3745 = w3717 ~^ in3[23];
assign w3746 = w2065 | w3718;
assign w3747 = w2267 | w3719;
assign w3748 = w2097 | w3720;
assign w3749 = w2173 | w3721;
assign w3750 = w1996 | w3722;
assign w3751 = w2324 | w3723;
assign w3752 = w2234 | w3724;
assign w3753 = w1187 | w3725;
assign w3754 = w1895 | w3726;
assign w3755 = w374 ~^ w3727;
assign w3756 = w375 | w3727;
assign w3757 = w3673 | w3731;
assign w3758 = w3676 | w3735;
assign w3759 = w3608 ~^ w3742;
assign w3760 = w3637 | w3742;
assign w3761 = ~w3742;
assign w3762 = ~w3744;
assign w3763 = w3612 ~^ w3745;
assign w3764 = w3639 | w3745;
assign w3765 = ~w3745;
assign w3766 = w2468 ~| w3746;
assign w3767 = w2592 ~| w3747;
assign w3768 = w2512 ~| w3748;
assign w3769 = w2543 ~| w3749;
assign w3770 = w2427 ~| w3750;
assign w3771 = w2627 ~| w3751;
assign w3772 = w2573 ~| w3752;
assign w3773 = w1152 ~| w3753;
assign w3774 = w2397 ~| w3754;
assign w3775 = w1245 ~| w3755;
assign w3776 = w1399 ~| w3755;
assign w3777 = w1295 ~| w3755;
assign w3778 = w837 ~| w3755;
assign w3779 = w1348 ~| w3755;
assign w3780 = w1486 ~| w3755;
assign w3781 = w1556 ~| w3755;
assign w3782 = w1522 ~| w3755;
assign w3783 = w1446 ~| w3755;
assign w3784 = w624 & w3756;
assign w3785 = w3736 ~^ w3759;
assign w3786 = w3736 & w3760;
assign w3787 = w3608 ~| w3761;
assign w3788 = w3732 ~^ w3763;
assign w3789 = w3732 & w3764;
assign w3790 = w3612 ~| w3765;
assign w3791 = w3766 ~^ in3[11];
assign w3792 = w3767 ~^ in3[23];
assign w3793 = w3768 ~^ in3[14];
assign w3794 = w3769 ~^ in3[17];
assign w3795 = w3770 ~^ in3[8];
assign w3796 = w3771 ~^ in3[26];
assign w3797 = w3772 ~^ in3[20];
assign w3798 = w3773 ~^ in3[2];
assign w3799 = w3774 ~^ in3[5];
assign w3800 = w1902 | w3775;
assign w3801 = w2085 | w3776;
assign w3802 = w1992 | w3777;
assign w3803 = w1194 | w3778;
assign w3804 = w2053 | w3779;
assign w3805 = w2248 | w3780;
assign w3806 = w2337 | w3781;
assign w3807 = w2262 | w3782;
assign w3808 = w2159 | w3783;
assign w3809 = w392 ~^ w3784;
assign w3810 = w393 | w3784;
assign w3811 = ~w3785;
assign w3812 = w3786 | w3787;
assign w3813 = ~w3788;
assign w3814 = w3789 | w3790;
assign w3815 = w3674 ~^ w3792;
assign w3816 = w3702 & w3792;
assign w3817 = w3669 ~^ w3796;
assign w3818 = w3700 & w3796;
assign w3819 = w2403 ~| w3800;
assign w3820 = w2522 ~| w3801;
assign w3821 = w2439 ~| w3802;
assign w3822 = w1157 ~| w3803;
assign w3823 = w2461 ~| w3804;
assign w3824 = w2564 ~| w3805;
assign w3825 = w2621 ~| w3806;
assign w3826 = w2611 ~| w3807;
assign w3827 = w2544 ~| w3808;
assign w3828 = w1291 ~| w3809;
assign w3829 = w831 ~| w3809;
assign w3830 = w1433 ~| w3809;
assign w3831 = w1482 ~| w3809;
assign w3832 = w1342 ~| w3809;
assign w3833 = w1524 ~| w3809;
assign w3834 = w1393 ~| w3809;
assign w3835 = w1239 ~| w3809;
assign w3836 = w625 & w3810;
assign w3837 = ~w3812;
assign w3838 = ~w3814;
assign w3839 = w3814 ~^ w3815;
assign w3840 = ~w3815;
assign w3841 = w3699 | w3816;
assign w3842 = w3812 ~^ w3817;
assign w3843 = ~w3817;
assign w3844 = w3698 | w3818;
assign w3845 = w3819 ~^ in3[5];
assign w3846 = w3820 ~^ in3[14];
assign w3847 = w3821 ~^ in3[8];
assign w3848 = w3822 ~^ in3[2];
assign w3849 = w3823 ~^ in3[11];
assign w3850 = w3824 ~^ in3[20];
assign w3851 = w3825 ~^ in3[26];
assign w3852 = w3826 ~^ in3[23];
assign w3853 = w3827 ~^ in3[17];
assign w3854 = w1999 | w3828;
assign w3855 = w1190 | w3829;
assign w3856 = w2193 | w3830;
assign w3857 = w2232 | w3831;
assign w3858 = w2008 | w3832;
assign w3859 = w2259 | w3833;
assign w3860 = w2072 | w3834;
assign w3861 = w1898 | w3835;
assign w3862 = w410 ~^ w3836;
assign w3863 = w411 | w3836;
assign w3864 = w3817 ~| w3837;
assign w3865 = w3815 ~| w3838;
assign w3866 = w3814 | w3840;
assign w3867 = ~w3841;
assign w3868 = w3812 | w3843;
assign w3869 = w3729 ~^ w3850;
assign w3870 = w3757 & w3850;
assign w3871 = w3728 ~^ w3851;
assign w3872 = w3733 ~^ w3852;
assign w3873 = w3758 & w3852;
assign w3874 = w2425 ~| w3854;
assign w3875 = w1139 ~| w3855;
assign w3876 = w2535 ~| w3856;
assign w3877 = w2578 ~| w3857;
assign w3878 = w2487 ~| w3858;
assign w3879 = w2606 ~| w3859;
assign w3880 = w2514 ~| w3860;
assign w3881 = w2407 ~| w3861;
assign w3882 = w1350 ~| w3862;
assign w3883 = w1518 ~| w3862;
assign w3884 = w1401 ~| w3862;
assign w3885 = w1247 ~| w3862;
assign w3886 = w1299 ~| w3862;
assign w3887 = w839 ~| w3862;
assign w3888 = w1447 ~| w3862;
assign w3889 = w1485 ~| w3862;
assign w3890 = w626 & w3863;
assign w3891 = ~w3869;
assign w3892 = w3730 | w3870;
assign w3893 = w3844 ~^ w3871;
assign w3894 = w3841 ~^ w3872;
assign w3895 = w3867 ~| w3872;
assign w3896 = ~w3872;
assign w3897 = w3734 | w3873;
assign w3898 = w3874 ~^ in3[8];
assign w3899 = w3875 ~^ in3[2];
assign w3900 = w3876 ~^ in3[17];
assign w3901 = w3877 ~^ in3[20];
assign w3902 = w3878 ~^ in3[11];
assign w3903 = w3879 ~^ in3[23];
assign w3904 = w3880 ~^ in3[14];
assign w3905 = w3881 ~^ in3[5];
assign w3906 = w2024 | w3882;
assign w3907 = w2271 | w3883;
assign w3908 = w2100 | w3884;
assign w3909 = w1904 | w3885;
assign w3910 = w2001 | w3886;
assign w3911 = w1196 | w3887;
assign w3912 = w2176 | w3888;
assign w3913 = w2224 | w3889;
assign w3914 = w428 ~^ w3890;
assign w3915 = w429 | w3890;
assign w3916 = w3841 | w3896;
assign w3917 = ~w3900;
assign w3918 = w3788 ~^ w3901;
assign w3919 = w3813 | w3901;
assign w3920 = ~w3901;
assign w3921 = w3785 ~^ w3903;
assign w3922 = w3811 | w3903;
assign w3923 = ~w3903;
assign w3924 = w2486 ~| w3906;
assign w3925 = w2596 ~| w3907;
assign w3926 = w2518 ~| w3908;
assign w3927 = w2413 ~| w3909;
assign w3928 = w2434 ~| w3910;
assign w3929 = w1135 ~| w3911;
assign w3930 = w2542 ~| w3912;
assign w3931 = w2559 ~| w3913;
assign w3932 = w838 ~| w3914;
assign w3933 = w1298 ~| w3914;
assign w3934 = w1246 ~| w3914;
assign w3935 = w1400 ~| w3914;
assign w3936 = w1519 ~| w3914;
assign w3937 = w1349 ~| w3914;
assign w3938 = w1490 ~| w3914;
assign w3939 = w1436 ~| w3914;
assign w3940 = w627 & w3915;
assign w3941 = w3892 ~^ w3918;
assign w3942 = w3892 & w3919;
assign w3943 = w3788 ~| w3920;
assign w3944 = w3897 ~^ w3921;
assign w3945 = w3897 & w3922;
assign w3946 = w3785 ~| w3923;
assign w3947 = w3924 ~^ in3[11];
assign w3948 = w3925 ~^ in3[23];
assign w3949 = w3926 ~^ in3[14];
assign w3950 = w3927 ~^ in3[5];
assign w3951 = w3928 ~^ in3[8];
assign w3952 = w3929 ~^ in3[2];
assign w3953 = w3930 ~^ in3[17];
assign w3954 = w3931 ~^ in3[20];
assign w3955 = w1175 | w3932;
assign w3956 = w1984 | w3933;
assign w3957 = w1883 | w3934;
assign w3958 = w2088 | w3935;
assign w3959 = w2261 | w3936;
assign w3960 = w2031 | w3937;
assign w3961 = w2231 | w3938;
assign w3962 = w2168 | w3939;
assign w3963 = w446 ~^ w3940;
assign w3964 = w447 | w3940;
assign w3965 = ~w3941;
assign w3966 = w3942 | w3943;
assign w3967 = ~w3944;
assign w3968 = w3945 | w3946;
assign w3969 = w3842 ~^ w3948;
assign w3970 = w3868 & w3948;
assign w3971 = w3839 ~^ w3954;
assign w3972 = w3866 & w3954;
assign w3973 = w1143 ~| w3955;
assign w3974 = w2441 ~| w3956;
assign w3975 = w2410 ~| w3957;
assign w3976 = w2508 ~| w3958;
assign w3977 = w2597 ~| w3959;
assign w3978 = w2481 ~| w3960;
assign w3979 = w2572 ~| w3961;
assign w3980 = w2540 ~| w3962;
assign w3981 = w1297 ~| w3963;
assign w3982 = w1484 ~| w3963;
assign w3983 = w835 ~| w3963;
assign w3984 = w1397 ~| w3963;
assign w3985 = w1445 ~| w3963;
assign w3986 = w1346 ~| w3963;
assign w3987 = w1243 ~| w3963;
assign w3988 = w628 & w3964;
assign w3989 = ~w3966;
assign w3990 = ~w3968;
assign w3991 = w3968 ~^ w3969;
assign w3992 = ~w3969;
assign w3993 = w3864 | w3970;
assign w3994 = w3966 ~^ w3971;
assign w3995 = ~w3971;
assign w3996 = w3865 | w3972;
assign w3997 = w3973 ~^ in3[2];
assign w3998 = w3974 ~^ in3[8];
assign w3999 = w3975 ~^ in3[5];
assign w4000 = w3976 ~^ in3[14];
assign w4001 = w3977 ~^ in3[23];
assign w4002 = w3978 ~^ in3[11];
assign w4003 = w3979 ~^ in3[20];
assign w4004 = w3980 ~^ in3[17];
assign w4005 = w2000 | w3981;
assign w4006 = w2242 | w3982;
assign w4007 = w1195 | w3983;
assign w4008 = w1367 | w3984;
assign w4009 = w2187 | w3985;
assign w4010 = w2027 | w3986;
assign w4011 = w1903 | w3987;
assign w4012 = w463 ~^ w3988;
assign w4013 = w464 | w3988;
assign w4014 = w3971 ~| w3989;
assign w4015 = w3969 ~| w3990;
assign w4016 = w3968 | w3992;
assign w4017 = w3966 | w3995;
assign w4018 = ~w3996;
assign w4019 = w3893 ~^ w4001;
assign w4020 = w3894 ~^ w4003;
assign w4021 = w3916 & w4003;
assign w4022 = w2436 ~| w4005;
assign w4023 = w2558 ~| w4006;
assign w4024 = w1164 ~| w4007;
assign w4025 = w2517 ~| w4008;
assign w4026 = w2534 ~| w4009;
assign w4027 = w2485 ~| w4010;
assign w4028 = w2415 ~| w4011;
assign w4029 = w823 ~| w4012;
assign w4030 = w1484 ~| w4012;
assign w4031 = w1283 ~| w4012;
assign w4032 = w1385 ~| w4012;
assign w4033 = w1444 ~| w4012;
assign w4034 = w1334 ~| w4012;
assign w4035 = w1233 ~| w4012;
assign w4036 = w629 & w4013;
assign w4037 = w3993 ~^ w4019;
assign w4038 = w3996 ~^ w4020;
assign w4039 = w4018 ~| w4020;
assign w4040 = ~w4020;
assign w4041 = w3895 | w4021;
assign w4042 = w4022 ~^ in3[8];
assign w4043 = w4023 ~^ in3[20];
assign w4044 = w4024 ~^ in3[2];
assign w4045 = w4025 ~^ in3[14];
assign w4046 = w4026 ~^ in3[17];
assign w4047 = w4027 ~^ in3[11];
assign w4048 = w4028 ~^ in3[5];
assign w4049 = w1189 | w4029;
assign w4050 = w2246 | w4030;
assign w4051 = w1964 | w4031;
assign w4052 = w2080 | w4032;
assign w4053 = w2171 | w4033;
assign w4054 = w2033 | w4034;
assign w4055 = w1897 | w4035;
assign w4056 = w479 ~^ w4036;
assign w4057 = w480 | w4036;
assign w4058 = w3996 | w4040;
assign w4059 = w3944 ~^ w4043;
assign w4060 = w3967 | w4043;
assign w4061 = ~w4043;
assign w4062 = ~w4045;
assign w4063 = w3941 ~^ w4046;
assign w4064 = w3965 | w4046;
assign w4065 = ~w4046;
assign w4066 = w1149 ~| w4049;
assign w4067 = w2567 ~| w4050;
assign w4068 = w2449 ~| w4051;
assign w4069 = w2513 ~| w4052;
assign w4070 = w2537 ~| w4053;
assign w4071 = w2483 ~| w4054;
assign w4072 = w2402 ~| w4055;
assign w4073 = w1388 ~| w4056;
assign w4074 = w1483 ~| w4056;
assign w4075 = w826 ~| w4056;
assign w4076 = w1337 ~| w4056;
assign w4077 = w1440 ~| w4056;
assign w4078 = w1286 ~| w4056;
assign w4079 = w1232 ~| w4056;
assign w4080 = w630 & w4057;
assign w4081 = w4041 ~^ w4059;
assign w4082 = w4041 & w4060;
assign w4083 = w3944 ~| w4061;
assign w4084 = w3941 ~| w4065;
assign w4085 = w4066 ~^ in3[2];
assign w4086 = w4067 ~^ in3[20];
assign w4087 = w4068 ~^ in3[8];
assign w4088 = w4069 ~^ in3[14];
assign w4089 = w4070 ~^ in3[17];
assign w4090 = w4071 ~^ in3[11];
assign w4091 = w4072 ~^ in3[5];
assign w4092 = w2093 | w4073;
assign w4093 = w2230 | w4074;
assign w4094 = w1193 | w4075;
assign w4095 = w2067 | w4076;
assign w4096 = w2178 | w4077;
assign w4097 = w1954 | w4078;
assign w4098 = w1901 | w4079;
assign w4099 = w494 ~^ w4080;
assign w4100 = w495 | w4080;
assign w4101 = ~w4081;
assign w4102 = w4082 | w4083;
assign w4103 = w3991 ~^ w4086;
assign w4104 = w4016 & w4086;
assign w4105 = w3994 ~^ w4089;
assign w4106 = w4017 & w4089;
assign w4107 = w2521 ~| w4092;
assign w4108 = w2563 ~| w4093;
assign w4109 = w1158 ~| w4094;
assign w4110 = w2465 ~| w4095;
assign w4111 = w2523 ~| w4096;
assign w4112 = w2451 ~| w4097;
assign w4113 = w2414 ~| w4098;
assign w4114 = w1284 ~| w4099;
assign w4115 = w1434 ~| w4099;
assign w4116 = w824 ~| w4099;
assign w4117 = w1335 ~| w4099;
assign w4118 = w1386 ~| w4099;
assign w4119 = w1234 ~| w4099;
assign w4120 = w631 & w4100;
assign w4121 = ~w4102;
assign w4122 = w4102 ~^ w4103;
assign w4123 = ~w4103;
assign w4124 = w4015 | w4104;
assign w4125 = ~w4105;
assign w4126 = w4014 | w4106;
assign w4127 = w4107 ~^ in3[14];
assign w4128 = w4108 ~^ in3[20];
assign w4129 = w4109 ~^ in3[2];
assign w4130 = w4110 ~^ in3[11];
assign w4131 = w4111 ~^ in3[17];
assign w4132 = w4112 ~^ in3[8];
assign w4133 = w4113 ~^ in3[5];
assign w4134 = w1963 | w4114;
assign w4135 = w2180 | w4115;
assign w4136 = w1182 | w4116;
assign w4137 = w2032 | w4117;
assign w4138 = w2087 | w4118;
assign w4139 = w1890 | w4119;
assign w4140 = w508 ~^ w4120;
assign w4141 = w509 | w4120;
assign w4142 = w4103 ~| w4121;
assign w4143 = w4102 | w4123;
assign w4144 = ~w4126;
assign w4145 = w4037 ~^ w4128;
assign w4146 = w4038 ~^ w4131;
assign w4147 = w4058 & w4131;
assign w4148 = w2446 ~| w4134;
assign w4149 = w2536 ~| w4135;
assign w4150 = w1159 ~| w4136;
assign w4151 = w2480 ~| w4137;
assign w4152 = w2511 ~| w4138;
assign w4153 = w2409 ~| w4139;
assign w4154 = w1396 ~| w4140;
assign w4155 = w1439 ~| w4140;
assign w4156 = w834 ~| w4140;
assign w4157 = w1296 ~| w4140;
assign w4158 = w1345 ~| w4140;
assign w4159 = w1242 ~| w4140;
assign w4160 = w632 & w4141;
assign w4161 = w4124 ~^ w4145;
assign w4162 = w4126 ~^ w4146;
assign w4163 = w4144 ~| w4146;
assign w4164 = ~w4146;
assign w4165 = w4039 | w4147;
assign w4166 = w4148 ~^ in3[8];
assign w4167 = w4149 ~^ in3[17];
assign w4168 = w4150 ~^ in3[2];
assign w4169 = w4151 ~^ in3[11];
assign w4170 = w4152 ~^ in3[14];
assign w4171 = w4153 ~^ in3[5];
assign w4172 = w2079 | w4154;
assign w4173 = w1419 | w4155;
assign w4174 = w1181 | w4156;
assign w4175 = w1961 | w4157;
assign w4176 = w2026 | w4158;
assign w4177 = w1889 | w4159;
assign w4178 = w519 ~^ w4160;
assign w4179 = w520 | w4160;
assign w4180 = w4126 | w4164;
assign w4181 = w4081 ~^ w4167;
assign w4182 = w4101 | w4167;
assign w4183 = ~w4167;
assign w4184 = ~w4169;
assign w4185 = ~w4170;
assign w4186 = w2510 ~| w4172;
assign w4187 = w2546 ~| w4173;
assign w4188 = w1165 ~| w4174;
assign w4189 = w2445 ~| w4175;
assign w4190 = w2479 ~| w4176;
assign w4191 = w2401 ~| w4177;
assign w4192 = w1340 ~| w4178;
assign w4193 = w1438 ~| w4178;
assign w4194 = w829 ~| w4178;
assign w4195 = w1391 ~| w4178;
assign w4196 = w1289 ~| w4178;
assign w4197 = w1237 ~| w4178;
assign w4198 = w633 & w4179;
assign w4199 = w4165 ~^ w4181;
assign w4200 = w4165 & w4182;
assign w4201 = w4081 ~| w4183;
assign w4202 = w4186 ~^ in3[14];
assign w4203 = w4187 ~^ in3[17];
assign w4204 = w4188 ~^ in3[2];
assign w4205 = w4189 ~^ in3[8];
assign w4206 = w4190 ~^ in3[11];
assign w4207 = w4191 ~^ in3[5];
assign w4208 = w2018 | w4192;
assign w4209 = w2170 | w4193;
assign w4210 = w1171 | w4194;
assign w4211 = w2099 | w4195;
assign w4212 = w1953 | w4196;
assign w4213 = w1933 | w4197;
assign w4214 = w530 ~^ w4198;
assign w4215 = w531 | w4198;
assign w4216 = ~w4199;
assign w4217 = w4200 | w4201;
assign w4218 = w4122 ~^ w4203;
assign w4219 = w4143 & w4203;
assign w4220 = w2475 ~| w4208;
assign w4221 = w2530 ~| w4209;
assign w4222 = w1155 ~| w4210;
assign w4223 = w2506 ~| w4211;
assign w4224 = w2443 ~| w4212;
assign w4225 = w2384 ~| w4213;
assign w4226 = w1297 ~| w4214;
assign w4227 = w835 ~| w4214;
assign w4228 = w1346 ~| w4214;
assign w4229 = w1397 ~| w4214;
assign w4230 = w1243 ~| w4214;
assign w4231 = w634 & w4215;
assign w4232 = ~w4217;
assign w4233 = w4217 ~^ w4218;
assign w4234 = ~w4218;
assign w4235 = w4142 | w4219;
assign w4236 = w4220 ~^ in3[11];
assign w4237 = w4221 ~^ in3[17];
assign w4238 = w4222 ~^ in3[2];
assign w4239 = w4223 ~^ in3[14];
assign w4240 = w4224 ~^ in3[8];
assign w4241 = w4225 ~^ in3[5];
assign w4242 = w1969 | w4226;
assign w4243 = w1167 | w4227;
assign w4244 = w2030 | w4228;
assign w4245 = w1352 | w4229;
assign w4246 = w1915 | w4230;
assign w4247 = w533 | w4231;
assign w4248 = ~w4231;
assign w4249 = w4218 ~| w4232;
assign w4250 = w4217 | w4234;
assign w4251 = w4161 ~^ w4237;
assign w4252 = w4162 ~^ w4239;
assign w4253 = w4180 & w4239;
assign w4254 = w2442 ~| w4242;
assign w4255 = w1150 ~| w4243;
assign w4256 = w2474 ~| w4244;
assign w4257 = w2504 ~| w4245;
assign w4258 = w2383 ~| w4246;
assign w4259 = w1390 ~| w4247;
assign w4260 = ~w4247;
assign w4261 = w828 ~| w4247;
assign w4262 = w1236 ~| w4247;
assign w4263 = w1288 ~| w4247;
assign w4264 = in1[31] ~| w4248;
assign w4265 = w4235 ~^ w4251;
assign w4266 = w4163 | w4253;
assign w4267 = w4254 ~^ in3[8];
assign w4268 = w4255 ~^ in3[2];
assign w4269 = w4256 ~^ in3[11];
assign w4270 = w4257 ~^ in3[14];
assign w4271 = w4258 ~^ in3[5];
assign w4272 = w2073 | w4259;
assign w4273 = ~w4260;
assign w4274 = w918 | w4261;
assign w4275 = w1907 | w4262;
assign w4276 = w1939 | w4263;
assign w4277 = w4260 | w4264;
assign w4278 = ~w4267;
assign w4279 = ~w4269;
assign w4280 = w4199 ~^ w4270;
assign w4281 = w4216 | w4270;
assign w4282 = ~w4270;
assign w4283 = w4272 ~^ in3[14];
assign w4284 = w1339 ~| w4273;
assign w4285 = w4274 ~^ in3[2];
assign w4286 = w4275 ~^ in3[5];
assign w4287 = w4276 ~^ in3[8];
assign w4288 = w1389 ~| w4277;
assign w4289 = w1338 ~| w4277;
assign w4290 = w1235 ~| w4277;
assign w4291 = w827 ~| w4277;
assign w4292 = w1287 ~| w4277;
assign w4293 = w4266 ~^ w4280;
assign w4294 = w4266 & w4281;
assign w4295 = w4199 ~| w4282;
assign w4296 = w4265 ~^ w4283;
assign w4297 = w2004 | w4284;
assign w4298 = ~w4286;
assign w4299 = ~w4287;
assign w4300 = w2488 ~| w4288;
assign w4301 = w2459 ~| w4289;
assign w4302 = w2392 ~| w4290;
assign w4303 = w1151 ~| w4291;
assign w4304 = w2421 ~| w4292;
assign w4305 = w4294 | w4295;
assign w4306 = w4297 ~^ in3[11];
assign w4307 = w4300 ~^ in3[14];
assign w4308 = w4301 ~^ in3[11];
assign w4309 = w4302 ~^ in3[5];
assign w4310 = w4303 ~^ in3[2];
assign w4311 = w4304 ~^ in3[8];
assign w4312 = ~w4305;
assign w4313 = ~w4306;
assign w4314 = w4233 ~^ w4307;
assign w4315 = w4250 & w4307;
assign w4316 = w4305 ~^ w4314;
assign w4317 = w4312 & w4314;
assign w4318 = w4312 ~| w4314;
assign w4319 = w4249 | w4315;
assign w4320 = w4296 ~^ w4319;
wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320;
endmodule
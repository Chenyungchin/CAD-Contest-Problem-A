module top(in1, in2, in3, out1);
input wire [18:0] in1;
input wire [18:0] in2;
input wire [18:0] in3;
output wire [19:0] out1;
assign w0 = ~in1[2];
assign w1 = ~in1[3];
assign w2 = ~in1[4];
assign w3 = ~in1[5];
assign w4 = ~in1[6];
assign w5 = ~in1[7];
assign w6 = ~in1[8];
assign w7 = ~in1[9];
assign w8 = ~in1[10];
assign w9 = ~in1[11];
assign w10 = ~in1[12];
assign w11 = ~in1[13];
assign w12 = ~in1[14];
assign w13 = ~in1[15];
assign w14 = ~in1[16];
assign w15 = ~in1[17];
assign w16 = in1[0] ~^ in2[0];
assign w17 = in1[0] & in2[0];
assign w18 = in1[0] | in2[0];
assign w19 = ~in2[1];
assign w20 = ~in2[2];
assign w21 = ~in2[3];
assign w22 = ~in2[4];
assign w23 = ~in2[5];
assign w24 = ~in2[7];
assign w25 = ~in2[8];
assign w26 = ~in2[9];
assign w27 = ~in2[10];
assign w28 = ~in2[11];
assign w29 = ~in2[12];
assign w30 = ~in2[13];
assign w31 = ~in2[14];
assign w32 = ~in2[15];
assign w33 = ~in2[16];
assign w34 = ~in2[17];
assign w35 = ~in2[18];
assign w36 = in3[1] & in2[1];
assign w37 = ~in3[1];
assign w38 = in3[2] ~^ in1[2];
assign w39 = ~in3[2];
assign w40 = in3[3] ~^ in1[3];
assign w41 = ~in3[3];
assign w42 = in3[4] ~^ in1[4];
assign w43 = ~in3[4];
assign w44 = in3[5] ~^ in1[5];
assign w45 = ~in3[5];
assign w46 = in3[6] ~^ in1[6];
assign w47 = ~in3[6];
assign w48 = in3[7] ~^ in1[7];
assign w49 = ~in3[7];
assign w50 = in3[8] ~^ in1[8];
assign w51 = ~in3[8];
assign w52 = in3[9] ~^ in1[9];
assign w53 = ~in3[9];
assign w54 = in3[10] ~^ in1[10];
assign w55 = ~in3[10];
assign w56 = in3[11] ~^ in1[11];
assign w57 = ~in3[11];
assign w58 = in3[12] ~^ in1[12];
assign w59 = ~in3[12];
assign w60 = in3[13] ~^ in1[13];
assign w61 = ~in3[13];
assign w62 = in3[14] ~^ in1[14];
assign w63 = ~in3[14];
assign w64 = in3[15] ~^ in1[15];
assign w65 = ~in3[15];
assign w66 = in3[16] ~^ in1[16];
assign w67 = ~in3[16];
assign w68 = in3[17] ~^ in1[17];
assign w69 = ~in3[17];
assign w70 = in3[18] ~^ in1[18];
assign w71 = in3[18] ~& in1[18];
assign out1[0] = w16 ~^ in3[0];
assign w72 = in3[0] & w18;
assign w73 = w19 & w37;
assign w74 = w20 | w38;
assign w75 = w20 & w38;
assign w76 = w0 | w39;
assign w77 = w40 ~^ in2[3];
assign w78 = w1 | w41;
assign w79 = w42 ~^ in2[4];
assign w80 = w2 | w43;
assign w81 = w3 & w45;
assign w82 = in2[6] ~| w46;
assign w83 = in2[6] & w46;
assign w84 = w4 & w47;
assign w85 = w48 ~^ in2[7];
assign w86 = w24 ~| w48;
assign w87 = w24 & w48;
assign w88 = w5 | w49;
assign w89 = w50 ~^ in2[8];
assign w90 = w25 & w50;
assign w91 = w25 ~| w50;
assign w92 = w6 | w51;
assign w93 = w52 ~^ in2[9];
assign w94 = w26 ~| w52;
assign w95 = w26 & w52;
assign w96 = w7 | w53;
assign w97 = w54 ~^ in2[10];
assign w98 = w8 | w55;
assign w99 = w56 ~^ in2[11];
assign w100 = w9 | w57;
assign w101 = w58 ~^ in2[12];
assign w102 = w10 | w59;
assign w103 = w60 ~^ in2[13];
assign w104 = w11 | w61;
assign w105 = w62 ~^ in2[14];
assign w106 = w12 | w63;
assign w107 = w64 ~^ in2[15];
assign w108 = w13 | w65;
assign w109 = w66 ~^ in2[16];
assign w110 = w14 | w67;
assign w111 = w68 ~^ in2[17];
assign w112 = w15 | w69;
assign w113 = w70 ~^ in2[18];
assign w114 = w35 & w70;
assign w115 = ~w70;
assign w116 = w17 | w72;
assign w117 = w36 | w73;
assign w118 = ~w75;
assign w119 = w21 & w76;
assign w120 = w21 ~| w76;
assign w121 = w76 ~^ w77;
assign w122 = w22 | w78;
assign w123 = ~w78;
assign w124 = w78 ~^ w79;
assign w125 = w80 ~^ in2[5];
assign w126 = w23 ~| w80;
assign w127 = ~w80;
assign w128 = w81 ~^ in2[6];
assign w129 = w81 ~| w82;
assign w130 = w84 ~^ w85;
assign w131 = w84 ~| w87;
assign w132 = w88 ~^ w89;
assign w133 = w88 ~| w90;
assign w134 = w92 ~^ w93;
assign w135 = w92 ~| w95;
assign w136 = w27 ~| w96;
assign w137 = w27 & w96;
assign w138 = w96 ~^ w97;
assign w139 = w28 ~| w98;
assign w140 = w28 & w98;
assign w141 = w98 ~^ w99;
assign w142 = w29 ~| w100;
assign w143 = w29 & w100;
assign w144 = w100 ~^ w101;
assign w145 = w30 ~| w102;
assign w146 = w30 & w102;
assign w147 = w102 ~^ w103;
assign w148 = w31 & w104;
assign w149 = w31 ~| w104;
assign w150 = w104 ~^ w105;
assign w151 = w32 ~| w106;
assign w152 = w32 & w106;
assign w153 = w106 ~^ w107;
assign w154 = w33 ~| w108;
assign w155 = w33 & w108;
assign w156 = w108 ~^ w109;
assign w157 = w34 ~| w110;
assign w158 = w34 & w110;
assign w159 = w110 ~^ w111;
assign w160 = w112 ~^ w113;
assign w161 = w112 ~| w114;
assign w162 = in2[18] & w115;
assign w163 = w117 ~^ in1[1];
assign w164 = in1[1] & w117;
assign w165 = in1[1] | w117;
assign w166 = w74 & w118;
assign w167 = w40 ~| w119;
assign w168 = w75 ~^ w121;
assign w169 = w118 ~| w121;
assign w170 = ~w121;
assign w171 = in2[4] ~| w123;
assign w172 = ~w124;
assign w173 = w44 ~^ w125;
assign w174 = in2[5] | w127;
assign w175 = w46 ~^ w128;
assign w176 = w83 | w129;
assign w177 = w86 | w131;
assign w178 = w91 | w133;
assign w179 = w94 | w135;
assign w180 = w54 ~| w137;
assign w181 = w56 ~| w140;
assign w182 = w58 ~| w143;
assign w183 = w60 ~| w146;
assign w184 = w62 ~| w148;
assign w185 = w64 ~| w152;
assign w186 = w66 ~| w155;
assign w187 = w68 ~| w158;
assign w188 = w161 ~| w162;
assign out1[1] = w116 ~^ w163;
assign w189 = w116 & w165;
assign w190 = w73 ~^ w166;
assign w191 = w73 | w166;
assign w192 = w73 & w166;
assign w193 = w120 | w167;
assign w194 = w75 | w170;
assign w195 = w42 | w171;
assign w196 = w44 & w174;
assign w197 = w130 ~^ w176;
assign w198 = w130 | w176;
assign w199 = w130 & w176;
assign w200 = w132 ~^ w177;
assign w201 = w132 & w177;
assign w202 = w132 | w177;
assign w203 = w134 ~^ w178;
assign w204 = w134 | w178;
assign w205 = w134 & w178;
assign w206 = w138 ~^ w179;
assign w207 = w138 | w179;
assign w208 = w138 & w179;
assign w209 = w136 | w180;
assign w210 = w139 | w181;
assign w211 = w142 | w182;
assign w212 = w145 | w183;
assign w213 = w149 | w184;
assign w214 = w151 | w185;
assign w215 = w154 | w186;
assign w216 = w157 | w187;
assign w217 = w71 ~^ w188;
assign w218 = w164 | w189;
assign w219 = w124 ~^ w193;
assign w220 = w124 ~| w193;
assign w221 = ~w193;
assign w222 = w122 & w195;
assign w223 = w126 | w196;
assign w224 = w141 ~^ w209;
assign w225 = w141 & w209;
assign w226 = w141 | w209;
assign w227 = w144 ~^ w210;
assign w228 = w144 & w210;
assign w229 = w144 | w210;
assign w230 = w147 ~^ w211;
assign w231 = w147 | w211;
assign w232 = w147 & w211;
assign w233 = w150 ~^ w212;
assign w234 = w150 & w212;
assign w235 = w150 | w212;
assign w236 = w153 ~^ w213;
assign w237 = w153 & w213;
assign w238 = w153 | w213;
assign w239 = w156 ~^ w214;
assign w240 = w156 | w214;
assign w241 = w156 & w214;
assign w242 = w159 ~^ w215;
assign w243 = w159 & w215;
assign w244 = w159 | w215;
assign w245 = w160 ~^ w216;
assign w246 = w160 & w216;
assign w247 = w160 | w216;
assign out1[2] = w190 ~^ w218;
assign w248 = ~w218;
assign w249 = w172 | w221;
assign w250 = w173 ~^ w222;
assign w251 = w173 | w222;
assign w252 = w173 & w222;
assign w253 = w175 ~^ w223;
assign w254 = ~w223;
assign w255 = w192 | w248;
assign w256 = w175 ~| w254;
assign w257 = w175 & w254;
assign w258 = w191 & w255;
assign out1[3] = w168 ~^ w258;
assign w259 = w169 | w258;
assign w260 = w194 & w259;
assign w261 = w220 | w260;
assign out1[4] = w219 ^ w260;
assign w262 = w249 & w261;
assign w263 = w252 | w262;
assign out1[5] = w250 ^ w262;
assign w264 = w251 & w263;
assign out1[6] = w253 ~^ w264;
assign w265 = w257 ~| w264;
assign w266 = w256 | w265;
assign out1[7] = w197 ~^ w266;
assign w267 = w198 & w266;
assign w268 = w199 | w267;
assign out1[8] = w200 ~^ w268;
assign w269 = w202 & w268;
assign w270 = w201 | w269;
assign out1[9] = w203 ~^ w270;
assign w271 = w204 & w270;
assign w272 = w205 | w271;
assign out1[10] = w206 ~^ w272;
assign w273 = w207 & w272;
assign w274 = w208 | w273;
assign out1[11] = w224 ~^ w274;
assign w275 = w226 & w274;
assign w276 = w225 | w275;
assign out1[12] = w227 ~^ w276;
assign w277 = w229 & w276;
assign w278 = w228 | w277;
assign out1[13] = w230 ~^ w278;
assign w279 = w231 & w278;
assign w280 = w232 | w279;
assign out1[14] = w233 ~^ w280;
assign w281 = w235 & w280;
assign w282 = w234 | w281;
assign out1[15] = w236 ~^ w282;
assign w283 = w238 & w282;
assign w284 = w237 | w283;
assign out1[16] = w239 ~^ w284;
assign w285 = w240 & w284;
assign w286 = w241 | w285;
assign out1[17] = w242 ~^ w286;
assign w287 = w244 & w286;
assign w288 = w243 | w287;
assign out1[18] = w245 ~^ w288;
assign w289 = w247 & w288;
assign w290 = w246 | w289;
assign out1[19] = w217 ~^ w290;
wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290;
endmodule
module top(in1, in2, in3, out1);
input wire [3:0] in1;
input wire [3:0] in2;
input wire [3:0] in3;
output wire [3:0] out1;
assign w0 = ~in1[0];
assign w1 = ~in1[1];
assign w2 = ~in1[2];
assign w3 = ~in1[3];
assign w4 = ~in2[0];
assign w5 = in1[1] & in2[1];
assign w6 = ~in2[1];
assign w7 = in1[0] & in2[2];
assign w8 = ~in2[2];
assign w9 = ~in2[3];
assign w10 = ~in3[0];
assign w11 = ~in3[2];
assign w12 = w1 | w4;
assign w13 = w2 | w4;
assign w14 = w0 | w4;
assign w15 = w3 | w4;
assign w16 = ~w5;
assign w17 = w2 | w6;
assign w18 = w0 | w6;
assign w19 = w5 | w7;
assign w20 = ~w7;
assign w21 = w1 | w8;
assign w22 = w0 | w9;
assign w23 = w12 ~^ in3[1];
assign w24 = ~w12;
assign w25 = w13 ~^ in3[2];
assign w26 = w11 | w13;
assign out1[0] = w14 ~^ in3[0];
assign w27 = w10 | w14;
assign w28 = w15 ~^ in3[3];
assign w29 = ~w18;
assign w30 = w16 ~^ w20;
assign w31 = w16 ~| w20;
assign w32 = w17 ~^ w22;
assign w33 = w18 ~^ w23;
assign w34 = ~w23;
assign w35 = in3[1] & w24;
assign w36 = w19 & w25;
assign w37 = w26 ~^ w28;
assign w38 = w23 ~| w29;
assign w39 = w25 ~^ w30;
assign w40 = w21 ~^ w32;
assign out1[1] = w27 ~^ w33;
assign w41 = w18 | w34;
assign w42 = w31 ~| w36;
assign w43 = w27 | w38;
assign w44 = w35 & w39;
assign w45 = w35 ~| w39;
assign w46 = w35 ^ w39;
assign w47 = w37 ~^ w40;
assign w48 = w41 & w43;
assign w49 = w42 ~^ w47;
assign out1[2] = w46 ~^ w48;
assign w50 = w45 ~| w48;
assign w51 = w44 ~| w50;
assign out1[3] = w49 ~^ w51;
wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51;
endmodule
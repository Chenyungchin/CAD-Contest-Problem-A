module top(in1, in2, in3, in4, out1);
input wire [15:0] in1;
input wire [15:0] in2;
input wire [15:0] in3;
input wire [1:0] in4;
output wire [31:0] out1;
assign w0 = ~in4[0];
assign w1 = in1[5] & in4[1];
assign w2 = in1[3] & in4[1];
assign w3 = in1[2] & in4[1];
assign w4 = in1[4] & in4[1];
assign w5 = in1[7] & in4[1];
assign w6 = in1[0] & in4[1];
assign w7 = in1[8] & in4[1];
assign w8 = in1[15] & in4[1];
assign w9 = in1[1] & in4[1];
assign w10 = in1[14] & in4[1];
assign w11 = in1[13] & in4[1];
assign w12 = in1[12] & in4[1];
assign w13 = in1[6] & in4[1];
assign w14 = in1[10] & in4[1];
assign w15 = in1[9] & in4[1];
assign w16 = in1[11] & in4[1];
assign w17 = in4[1] | in4[0];
assign w18 = ~in4[1];
assign w19 = ~in4[1];
assign w20 = ~in4[1];
assign w21 = ~in4[1];
assign w22 = ~in4[1];
assign w23 = ~in4[1];
assign w24 = ~in4[1];
assign w25 = ~in4[1];
assign w26 = ~in4[1];
assign w27 = in2[4] & w18;
assign w28 = in2[6] & w18;
assign w29 = w0 | w18;
assign w30 = in2[2] & w19;
assign w31 = in2[10] & w19;
assign w32 = in2[8] & w20;
assign w33 = in2[0] & w21;
assign w34 = in2[12] & w21;
assign w35 = in2[3] & w22;
assign w36 = in2[11] & w22;
assign w37 = in2[15] & w23;
assign w38 = in2[14] & w23;
assign w39 = in2[7] & w24;
assign w40 = in2[5] & w25;
assign w41 = in2[13] & w25;
assign w42 = in2[1] & w26;
assign w43 = in2[9] & w26;
assign w44 = w4 | w27;
assign w45 = w13 | w28;
assign w46 = w17 & w29;
assign w47 = ~w29;
assign w48 = ~w29;
assign w49 = ~w29;
assign w50 = ~w29;
assign w51 = ~w29;
assign w52 = ~w29;
assign w53 = ~w29;
assign w54 = ~w29;
assign w55 = w3 | w30;
assign w56 = w14 | w31;
assign w57 = w7 | w32;
assign w58 = w6 | w33;
assign w59 = w12 | w34;
assign w60 = w2 | w35;
assign w61 = w16 | w36;
assign w62 = w8 | w37;
assign w63 = w10 | w38;
assign w64 = w5 | w39;
assign w65 = w1 | w40;
assign w66 = w11 | w41;
assign w67 = w9 | w42;
assign w68 = w15 | w43;
assign w69 = ~w44;
assign w70 = ~w45;
assign w71 = in3[3] & w46;
assign w72 = in3[1] & w46;
assign w73 = in3[0] & w46;
assign w74 = in3[9] & w46;
assign w75 = in3[10] & w46;
assign w76 = in3[7] & w46;
assign w77 = in3[14] & w46;
assign w78 = in3[8] & w46;
assign w79 = in3[12] & w46;
assign w80 = in3[6] & w46;
assign w81 = in3[4] & w46;
assign w82 = in3[11] & w46;
assign w83 = in3[2] & w46;
assign w84 = in3[5] & w46;
assign w85 = in3[13] & w46;
assign w86 = in3[15] & w46;
assign w87 = in2[3] & w47;
assign w88 = in2[8] & w47;
assign w89 = in2[15] & w48;
assign w90 = in2[11] & w48;
assign w91 = in2[1] & w49;
assign w92 = in2[4] & w49;
assign w93 = in2[12] & w50;
assign w94 = in2[5] & w50;
assign w95 = in2[10] & w51;
assign w96 = in2[7] & w51;
assign w97 = in2[2] & w52;
assign w98 = in2[9] & w52;
assign w99 = in2[13] & w53;
assign w100 = in2[14] & w53;
assign w101 = in2[0] & w54;
assign w102 = in2[6] & w54;
assign w103 = ~w55;
assign w104 = ~w55;
assign w105 = ~w55;
assign w106 = ~w55;
assign w107 = ~w56;
assign w108 = ~w57;
assign w109 = ~w57;
assign w110 = ~w57;
assign w111 = ~w57;
assign w112 = ~w57;
assign w113 = ~w57;
assign w114 = ~w57;
assign w115 = ~w57;
assign w116 = ~w57;
assign w117 = ~w57;
assign w118 = ~w58;
assign w119 = ~w59;
assign w120 = ~w60;
assign w121 = w55 ~^ w60;
assign w122 = ~w61;
assign w123 = ~w61;
assign w124 = ~w61;
assign w125 = ~w61;
assign w126 = ~w61;
assign w127 = ~w61;
assign w128 = ~w61;
assign w129 = ~w61;
assign w130 = ~w61;
assign w131 = ~w61;
assign w132 = ~w62;
assign w133 = ~w63;
assign w134 = ~w63;
assign w135 = ~w63;
assign w136 = ~w63;
assign w137 = ~w63;
assign w138 = ~w63;
assign w139 = w62 | w63;
assign w140 = ~w63;
assign w141 = ~w63;
assign w142 = ~w64;
assign w143 = ~w65;
assign w144 = ~w65;
assign w145 = ~w65;
assign w146 = ~w65;
assign w147 = ~w65;
assign w148 = w55 ~| w65;
assign w149 = ~w65;
assign w150 = ~w65;
assign w151 = ~w65;
assign w152 = ~w65;
assign w153 = ~w66;
assign w154 = ~w67;
assign w155 = ~w68;
assign w156 = w60 | w69;
assign w157 = ~w69;
assign w158 = w64 | w70;
assign w159 = w71 | w87;
assign w160 = w78 | w88;
assign w161 = w86 | w89;
assign w162 = w82 | w90;
assign w163 = w72 | w91;
assign w164 = w81 | w92;
assign w165 = w79 | w93;
assign w166 = w84 | w94;
assign w167 = w75 | w95;
assign w168 = w76 | w96;
assign w169 = w83 | w97;
assign w170 = w74 | w98;
assign w171 = w85 | w99;
assign w172 = w77 | w100;
assign w173 = w73 | w101;
assign w174 = w80 | w102;
assign w175 = w67 | w105;
assign w176 = w67 ~^ w105;
assign w177 = ~w106;
assign w178 = w68 | w107;
assign w179 = ~w108;
assign w180 = ~w109;
assign w181 = ~w110;
assign w182 = ~w111;
assign w183 = ~w112;
assign w184 = ~w113;
assign w185 = w66 | w119;
assign w186 = ~w122;
assign w187 = ~w123;
assign w188 = ~w124;
assign w189 = ~w125;
assign w190 = ~w126;
assign w191 = ~w127;
assign w192 = ~w128;
assign w193 = w119 ~^ w131;
assign w194 = ~w133;
assign w195 = ~w134;
assign w196 = ~w135;
assign w197 = ~w136;
assign w198 = ~w137;
assign w199 = ~w138;
assign w200 = w132 | w140;
assign w201 = w45 | w142;
assign w202 = ~w143;
assign w203 = ~w144;
assign w204 = ~w145;
assign w205 = ~w146;
assign w206 = ~w147;
assign w207 = w44 ~^ w150;
assign w208 = w105 | w151;
assign w209 = w55 & w151;
assign w210 = w70 ~^ w152;
assign w211 = w59 | w153;
assign w212 = w58 | w154;
assign w213 = w116 ~^ w155;
assign w214 = w56 | w155;
assign w215 = w55 | w156;
assign w216 = w120 | w157;
assign w217 = w149 | w158;
assign w218 = ~w159;
assign w219 = ~w159;
assign w220 = ~w159;
assign w221 = ~w159;
assign w222 = ~w159;
assign w223 = ~w159;
assign w224 = ~w159;
assign w225 = ~w159;
assign w226 = ~w159;
assign w227 = ~w159;
assign w228 = ~w160;
assign w229 = ~w160;
assign w230 = ~w160;
assign w231 = ~w160;
assign w232 = ~w160;
assign w233 = ~w160;
assign w234 = ~w160;
assign w235 = ~w160;
assign w236 = ~w160;
assign w237 = ~w160;
assign w238 = ~w161;
assign w239 = ~w161;
assign w240 = ~w161;
assign w241 = ~w161;
assign w242 = ~w161;
assign w243 = ~w161;
assign w244 = ~w161;
assign w245 = ~w161;
assign w246 = ~w161;
assign w247 = ~w161;
assign w248 = ~w162;
assign w249 = ~w162;
assign w250 = ~w162;
assign w251 = ~w162;
assign w252 = ~w162;
assign w253 = ~w162;
assign w254 = ~w162;
assign w255 = ~w162;
assign w256 = ~w162;
assign w257 = ~w162;
assign w258 = ~w163;
assign w259 = ~w163;
assign w260 = ~w163;
assign w261 = ~w163;
assign w262 = ~w163;
assign w263 = ~w163;
assign w264 = ~w163;
assign w265 = ~w163;
assign w266 = w159 ~| w164;
assign w267 = w159 ~^ w164;
assign w268 = ~w164;
assign w269 = ~w164;
assign w270 = ~w164;
assign w271 = ~w164;
assign w272 = ~w164;
assign w273 = ~w164;
assign w274 = ~w164;
assign w275 = ~w164;
assign w276 = ~w164;
assign w277 = ~w164;
assign w278 = w162 ~^ w165;
assign w279 = w162 ~| w165;
assign w280 = ~w165;
assign w281 = ~w165;
assign w282 = ~w165;
assign w283 = ~w165;
assign w284 = ~w165;
assign w285 = ~w165;
assign w286 = ~w165;
assign w287 = ~w165;
assign w288 = ~w165;
assign w289 = ~w165;
assign w290 = w164 ~^ w166;
assign w291 = w164 ~| w166;
assign w292 = ~w166;
assign w293 = ~w166;
assign w294 = ~w166;
assign w295 = ~w166;
assign w296 = ~w166;
assign w297 = ~w166;
assign w298 = ~w166;
assign w299 = ~w166;
assign w300 = ~w166;
assign w301 = ~w166;
assign w302 = w162 ~^ w167;
assign w303 = w162 ~| w167;
assign w304 = ~w167;
assign w305 = ~w167;
assign w306 = ~w167;
assign w307 = ~w167;
assign w308 = ~w167;
assign w309 = ~w167;
assign w310 = ~w167;
assign w311 = ~w167;
assign w312 = ~w167;
assign w313 = ~w167;
assign w314 = w160 ~| w168;
assign w315 = w160 ~^ w168;
assign w316 = ~w168;
assign w317 = ~w168;
assign w318 = ~w168;
assign w319 = ~w168;
assign w320 = ~w168;
assign w321 = ~w168;
assign w322 = ~w168;
assign w323 = ~w168;
assign w324 = ~w168;
assign w325 = ~w168;
assign w326 = w159 ~| w169;
assign w327 = w163 ~^ w169;
assign w328 = w159 ~^ w169;
assign w329 = ~w169;
assign w330 = ~w169;
assign w331 = ~w169;
assign w332 = ~w169;
assign w333 = ~w169;
assign w334 = ~w169;
assign w335 = ~w169;
assign w336 = ~w169;
assign w337 = ~w169;
assign w338 = ~w169;
assign w339 = w160 ~| w170;
assign w340 = w167 ~| w170;
assign w341 = w160 ~^ w170;
assign w342 = w167 ~^ w170;
assign w343 = ~w170;
assign w344 = ~w170;
assign w345 = ~w170;
assign w346 = ~w170;
assign w347 = ~w170;
assign w348 = ~w170;
assign w349 = ~w170;
assign w350 = ~w170;
assign w351 = ~w170;
assign w352 = ~w170;
assign w353 = w165 ~| w171;
assign w354 = w165 ~^ w171;
assign w355 = ~w171;
assign w356 = ~w171;
assign w357 = ~w171;
assign w358 = ~w171;
assign w359 = ~w171;
assign w360 = ~w171;
assign w361 = ~w171;
assign w362 = ~w171;
assign w363 = ~w171;
assign w364 = ~w171;
assign w365 = w171 ~| w172;
assign w366 = w161 ~| w172;
assign w367 = w171 ~^ w172;
assign w368 = w161 ~^ w172;
assign w369 = ~w172;
assign w370 = ~w172;
assign w371 = ~w172;
assign w372 = ~w172;
assign w373 = ~w172;
assign w374 = ~w172;
assign w375 = ~w172;
assign w376 = ~w172;
assign w377 = ~w172;
assign w378 = ~w172;
assign w379 = w163 ~^ w173;
assign w380 = ~w173;
assign w381 = ~w173;
assign w382 = ~w173;
assign w383 = ~w173;
assign w384 = ~w173;
assign w385 = w168 ~| w174;
assign w386 = w166 ~| w174;
assign w387 = w166 ~^ w174;
assign w388 = w168 ~^ w174;
assign w389 = ~w174;
assign w390 = ~w174;
assign w391 = ~w174;
assign w392 = ~w174;
assign w393 = ~w174;
assign w394 = ~w174;
assign w395 = ~w174;
assign w396 = ~w174;
assign w397 = ~w174;
assign w398 = ~w174;
assign w399 = w58 | w175;
assign w400 = w118 | w176;
assign w401 = ~w176;
assign w402 = w142 | w180;
assign w403 = w178 | w181;
assign w404 = w142 & w183;
assign w405 = w130 | w185;
assign w406 = w107 & w187;
assign w407 = w107 | w192;
assign w408 = w153 | w194;
assign w409 = w153 & w197;
assign w410 = w139 & w200;
assign w411 = w105 & w203;
assign w412 = w201 | w204;
assign w413 = w121 | w207;
assign w414 = ~w207;
assign w415 = w44 & w209;
assign w416 = w190 | w211;
assign w417 = w116 | w214;
assign w418 = w103 | w216;
assign w419 = w200 ~| w219;
assign w420 = w212 ~| w224;
assign w421 = w212 ~| w229;
assign w422 = w200 ~| w234;
assign w423 = w212 ~| w239;
assign w424 = w200 | w239;
assign w425 = w212 ~| w249;
assign w426 = w200 ~| w254;
assign w427 = w200 ~| w258;
assign w428 = w212 ~| w262;
assign w429 = w200 ~| w269;
assign w430 = w212 ~| w274;
assign w431 = w224 | w274;
assign w432 = w200 ~| w281;
assign w433 = w212 ~| w286;
assign w434 = w249 | w286;
assign w435 = w200 ~| w293;
assign w436 = w212 ~| w298;
assign w437 = w269 | w298;
assign w438 = w212 ~| w305;
assign w439 = w254 | w305;
assign w440 = w200 ~| w310;
assign w441 = w200 ~| w317;
assign w442 = w229 | w317;
assign w443 = w212 ~| w322;
assign w444 = w200 ~| w330;
assign w445 = w219 | w330;
assign w446 = w212 ~| w335;
assign w447 = w258 | w335;
assign w448 = w212 ~| w344;
assign w449 = w310 | w344;
assign w450 = w200 ~| w349;
assign w451 = w234 | w349;
assign w452 = w212 ~| w356;
assign w453 = w281 | w356;
assign w454 = w200 ~| w361;
assign w455 = w212 ~| w370;
assign w456 = w247 | w370;
assign w457 = w200 ~| w375;
assign w458 = w361 | w375;
assign w459 = w212 ~| w382;
assign w460 = w200 ~| w383;
assign w461 = w262 | w384;
assign w462 = w200 ~| w390;
assign w463 = w293 | w390;
assign w464 = w212 ~| w395;
assign w465 = w322 | w395;
assign w466 = w295 ~| w399;
assign w467 = w381 ~| w399;
assign w468 = w283 ~| w399;
assign w469 = w358 ~| w399;
assign w470 = w221 ~| w399;
assign w471 = w271 ~| w399;
assign w472 = w372 ~| w399;
assign w473 = w332 ~| w399;
assign w474 = w307 ~| w399;
assign w475 = w251 ~| w399;
assign w476 = w260 ~| w399;
assign w477 = w231 ~| w399;
assign w478 = w319 ~| w399;
assign w479 = w346 ~| w399;
assign w480 = w392 ~| w399;
assign w481 = w244 ~| w399;
assign w482 = w262 ~| w400;
assign w483 = w284 ~| w400;
assign w484 = w318 ~| w400;
assign w485 = w272 ~| w400;
assign w486 = w360 ~| w400;
assign w487 = w369 ~| w400;
assign w488 = w334 ~| w400;
assign w489 = w312 ~| w400;
assign w490 = w240 ~| w400;
assign w491 = w389 ~| w400;
assign w492 = w292 ~| w400;
assign w493 = w226 ~| w400;
assign w494 = w345 ~| w400;
assign w495 = w256 ~| w400;
assign w496 = w230 ~| w400;
assign w497 = w118 | w401;
assign w498 = w70 | w402;
assign w499 = ~w402;
assign w500 = ~w404;
assign w501 = ~w406;
assign w502 = w155 | w407;
assign w503 = ~w407;
assign w504 = w119 | w408;
assign w505 = ~w408;
assign w506 = ~w409;
assign w507 = w173 & w410;
assign w508 = w166 & w410;
assign w509 = w163 & w410;
assign w510 = w169 & w410;
assign w511 = w160 & w410;
assign w512 = w174 & w410;
assign w513 = w168 & w410;
assign w514 = w172 & w410;
assign w515 = w161 & w410;
assign w516 = w162 & w410;
assign w517 = w167 & w410;
assign w518 = w164 & w410;
assign w519 = w171 & w410;
assign w520 = w159 & w410;
assign w521 = w170 & w410;
assign w522 = w165 & w410;
assign w523 = w209 ~| w411;
assign w524 = ~w411;
assign w525 = w217 & w412;
assign w526 = w220 ~| w413;
assign w527 = w393 ~| w413;
assign w528 = w320 ~| w413;
assign w529 = w363 ~| w413;
assign w530 = w242 ~| w413;
assign w531 = w347 ~| w413;
assign w532 = w306 ~| w413;
assign w533 = w250 ~| w413;
assign w534 = w263 ~| w413;
assign w535 = w300 ~| w413;
assign w536 = w228 ~| w413;
assign w537 = w268 ~| w413;
assign w538 = w331 ~| w413;
assign w539 = w374 ~| w413;
assign w540 = w282 ~| w413;
assign w541 = w121 | w414;
assign w542 = w60 & w415;
assign w543 = w405 & w416;
assign w544 = w403 & w417;
assign w545 = w215 & w418;
assign w546 = w447 & w461;
assign w547 = w464 | w466;
assign w548 = w428 | w467;
assign w549 = w452 | w468;
assign w550 = w455 | w469;
assign w551 = w430 | w470;
assign w552 = w436 | w471;
assign w553 = w423 | w472;
assign w554 = w420 | w473;
assign w555 = w425 | w474;
assign w556 = w433 | w475;
assign w557 = w446 | w476;
assign w558 = w448 | w477;
assign w559 = w421 | w478;
assign w560 = w438 | w479;
assign w561 = w443 | w480;
assign w562 = w459 | w482;
assign w563 = w400 & w497;
assign w564 = w379 ~| w497;
assign w565 = w149 ~| w498;
assign w566 = w404 | w499;
assign w567 = w45 ~| w500;
assign w568 = w68 ~| w501;
assign w569 = w114 ~| w502;
assign w570 = w406 | w503;
assign w571 = w129 ~| w504;
assign w572 = w409 | w505;
assign w573 = w59 ~| w506;
assign w574 = ~w507;
assign w575 = w429 | w508;
assign w576 = w460 | w509;
assign w577 = w427 | w510;
assign w578 = w441 | w511;
assign w579 = w435 | w512;
assign w580 = w462 | w513;
assign w581 = w454 | w514;
assign w582 = w457 | w515;
assign w583 = w440 | w516;
assign w584 = w450 | w517;
assign w585 = w419 | w518;
assign w586 = w432 | w519;
assign w587 = w444 | w520;
assign w588 = w422 | w521;
assign w589 = w426 | w522;
assign w590 = w157 | w524;
assign w591 = w380 ~| w525;
assign w592 = w222 ~| w525;
assign w593 = w232 ~| w525;
assign w594 = w329 ~| w525;
assign w595 = w258 ~| w525;
assign w596 = w321 ~| w525;
assign w597 = w373 ~| w525;
assign w598 = w355 ~| w525;
assign w599 = w241 ~| w525;
assign w600 = w351 ~| w525;
assign w601 = w297 ~| w525;
assign w602 = w394 ~| w525;
assign w603 = w308 ~| w525;
assign w604 = w288 ~| w525;
assign w605 = w253 ~| w525;
assign w606 = w272 ~| w525;
assign w607 = w413 & w541;
assign w608 = w379 ~| w541;
assign w609 = w382 ~| w543;
assign w610 = w359 ~| w543;
assign w611 = w244 ~| w543;
assign w612 = w333 ~| w543;
assign w613 = w252 ~| w543;
assign w614 = w285 ~| w543;
assign w615 = w371 ~| w543;
assign w616 = w348 ~| w543;
assign w617 = w261 ~| w543;
assign w618 = w218 ~| w543;
assign w619 = w324 ~| w543;
assign w620 = w273 ~| w543;
assign w621 = w294 ~| w543;
assign w622 = w308 ~| w543;
assign w623 = w232 ~| w543;
assign w624 = w397 ~| w543;
assign w625 = w381 ~| w544;
assign w626 = w222 ~| w544;
assign w627 = w309 ~| w544;
assign w628 = w343 ~| w544;
assign w629 = w284 ~| w544;
assign w630 = w233 ~| w544;
assign w631 = w296 ~| w544;
assign w632 = w276 ~| w544;
assign w633 = w264 ~| w544;
assign w634 = w252 ~| w544;
assign w635 = w243 ~| w544;
assign w636 = w373 ~| w544;
assign w637 = w359 ~| w544;
assign w638 = w333 ~| w544;
assign w639 = w316 ~| w544;
assign w640 = w391 ~| w544;
assign w641 = w380 ~| w545;
assign w642 = w296 ~| w545;
assign w643 = w270 ~| w545;
assign w644 = w337 ~| w545;
assign w645 = w347 ~| w545;
assign w646 = w393 ~| w545;
assign w647 = w280 ~| w545;
assign w648 = w223 ~| w545;
assign w649 = w261 ~| w545;
assign w650 = w236 ~| w545;
assign w651 = w377 ~| w545;
assign w652 = w304 ~| w545;
assign w653 = w320 ~| w545;
assign w654 = w248 ~| w545;
assign w655 = w357 ~| w545;
assign w656 = w241 ~| w545;
assign w657 = w328 ~^ w546;
assign w658 = w326 | w546;
assign w659 = w381 | w563;
assign w660 = w562 ~| w564;
assign w661 = w210 | w566;
assign w662 = ~w566;
assign w663 = w150 & w567;
assign w664 = w117 & w568;
assign w665 = w213 | w570;
assign w666 = ~w570;
assign w667 = w193 | w572;
assign w668 = ~w572;
assign w669 = w131 & w573;
assign w670 = w55 ~^ w575;
assign w671 = w55 | w575;
assign w672 = w55 & w575;
assign w673 = ~w578;
assign w674 = w115 & w578;
assign w675 = w523 ~^ w579;
assign w676 = w208 & w579;
assign w677 = ~w580;
assign w678 = ~w581;
assign w679 = w133 ^ w582;
assign w680 = ~w583;
assign w681 = w130 | w583;
assign w682 = ~w584;
assign w683 = w55 ~^ w585;
assign w684 = w55 & w585;
assign w685 = w55 | w585;
assign w686 = w581 ~^ w586;
assign w687 = w140 | w586;
assign w688 = w55 ~^ w587;
assign w689 = w55 & w587;
assign w690 = w55 | w587;
assign w691 = w111 ^ w588;
assign w692 = w122 ^ w589;
assign w693 = w60 ~| w590;
assign w694 = w384 | w607;
assign w695 = w534 | w641;
assign w696 = w527 | w642;
assign w697 = w532 | w645;
assign w698 = w528 | w646;
assign w699 = w538 | w649;
assign w700 = w531 | w650;
assign w701 = w530 | w651;
assign w702 = w533 | w652;
assign w703 = w536 | w653;
assign w704 = w541 ~| w657;
assign w705 = w497 ~| w657;
assign w706 = w445 & w658;
assign w707 = w105 ^ w659;
assign w708 = w104 ~^ w660;
assign w709 = w260 ~| w661;
assign w710 = w256 ~| w661;
assign w711 = w324 ~| w661;
assign w712 = w312 ~| w661;
assign w713 = w295 ~| w661;
assign w714 = w358 ~| w661;
assign w715 = w276 ~| w661;
assign w716 = w376 ~| w661;
assign w717 = w242 ~| w661;
assign w718 = w350 ~| w661;
assign w719 = w235 ~| w661;
assign w720 = w225 ~| w661;
assign w721 = w396 ~| w661;
assign w722 = w336 ~| w661;
assign w723 = w288 ~| w661;
assign w724 = w210 | w662;
assign w725 = w565 | w663;
assign w726 = w569 | w664;
assign w727 = w351 ~| w665;
assign w728 = w300 ~| w665;
assign w729 = w238 ~| w665;
assign w730 = w264 ~| w665;
assign w731 = w323 ~| w665;
assign w732 = w251 ~| w665;
assign w733 = w377 ~| w665;
assign w734 = w231 ~| w665;
assign w735 = w397 ~| w665;
assign w736 = w275 ~| w665;
assign w737 = w311 ~| w665;
assign w738 = w287 ~| w665;
assign w739 = w363 ~| w665;
assign w740 = w226 ~| w665;
assign w741 = w332 ~| w665;
assign w742 = w213 | w666;
assign w743 = w337 ~| w667;
assign w744 = w319 ~| w667;
assign w745 = w259 ~| w667;
assign w746 = w307 ~| w667;
assign w747 = w283 ~| w667;
assign w748 = w255 ~| w667;
assign w749 = w362 ~| w667;
assign w750 = w236 ~| w667;
assign w751 = w392 ~| w667;
assign w752 = w221 ~| w667;
assign w753 = w372 ~| w667;
assign w754 = w299 ~| w667;
assign w755 = w245 ~| w667;
assign w756 = w271 ~| w667;
assign w757 = w346 ~| w667;
assign w758 = w193 | w668;
assign w759 = w571 | w669;
assign w760 = w580 | w673;
assign w761 = ~w673;
assign w762 = w148 | w676;
assign w763 = w578 ~| w677;
assign w764 = w586 | w678;
assign w765 = w584 | w680;
assign w766 = ~w680;
assign w767 = w589 & w681;
assign w768 = w583 ~| w682;
assign w769 = w582 & w687;
assign w770 = w578 ~^ w691;
assign w771 = w583 ~^ w692;
assign w772 = w542 | w693;
assign w773 = w65 ~^ w694;
assign w774 = w608 ~| w695;
assign w775 = w526 | w704;
assign w776 = w493 | w705;
assign w777 = w267 ~^ w706;
assign w778 = w266 | w706;
assign out1[0] = w104 ~^ w707;
assign w779 = ~w707;
assign w780 = w604 | w714;
assign w781 = w595 | w722;
assign w782 = w605 | w723;
assign w783 = w657 ~| w724;
assign w784 = w661 & w724;
assign w785 = w379 ~| w724;
assign w786 = ~w725;
assign w787 = ~w725;
assign w788 = ~w725;
assign w789 = ~w725;
assign w790 = ~w725;
assign w791 = w173 & w725;
assign w792 = ~w725;
assign w793 = ~w725;
assign w794 = ~w726;
assign w795 = ~w726;
assign w796 = ~w726;
assign w797 = ~w726;
assign w798 = ~w726;
assign w799 = w173 & w726;
assign w800 = ~w726;
assign w801 = ~w726;
assign w802 = w632 | w728;
assign w803 = w625 | w730;
assign w804 = w626 | w736;
assign w805 = w628 | w737;
assign w806 = w638 | w740;
assign w807 = w633 | w741;
assign w808 = ~w742;
assign w809 = w379 ~| w742;
assign w810 = w617 | w743;
assign w811 = w624 | w744;
assign w812 = w609 | w745;
assign w813 = w621 | w751;
assign w814 = w612 | w752;
assign w815 = w620 | w754;
assign w816 = w618 | w756;
assign w817 = w657 ~| w758;
assign w818 = w667 & w758;
assign w819 = w379 ~| w758;
assign w820 = ~w759;
assign w821 = ~w759;
assign w822 = ~w759;
assign w823 = ~w759;
assign w824 = ~w759;
assign w825 = w173 & w759;
assign w826 = ~w759;
assign w827 = ~w759;
assign w828 = w580 ~^ w761;
assign w829 = w115 | w761;
assign w830 = w580 ~^ w762;
assign w831 = w677 | w762;
assign w832 = w677 & w762;
assign w833 = w584 ~^ w766;
assign w834 = w129 & w766;
assign w835 = ~w770;
assign w836 = ~w771;
assign w837 = ~w772;
assign w838 = ~w772;
assign w839 = ~w772;
assign w840 = ~w772;
assign w841 = ~w772;
assign w842 = w173 & w772;
assign w843 = ~w772;
assign w844 = ~w772;
assign w845 = ~w773;
assign w846 = w143 ^ w773;
assign w847 = w206 ~^ w774;
assign w848 = w557 ~| w776;
assign w849 = w724 ~| w777;
assign w850 = w742 ~| w777;
assign w851 = w497 ~| w777;
assign w852 = w758 ~| w777;
assign w853 = w541 ~| w777;
assign w854 = w431 & w778;
assign w855 = w103 | w779;
assign w856 = w720 | w783;
assign w857 = w382 | w784;
assign w858 = w591 | w785;
assign w859 = w227 ~| w786;
assign w860 = w273 ~| w786;
assign w861 = w285 ~| w786;
assign w862 = w238 ~| w787;
assign w863 = w316 ~| w787;
assign w864 = w259 ~| w788;
assign w865 = w355 ~| w788;
assign w866 = w338 ~| w789;
assign w867 = w398 ~| w789;
assign w868 = w257 ~| w790;
assign w869 = w237 ~| w790;
assign w870 = w352 ~| w792;
assign w871 = w297 ~| w792;
assign w872 = w313 ~| w793;
assign w873 = w369 ~| w793;
assign w874 = w329 ~| w794;
assign w875 = w374 ~| w794;
assign w876 = w248 ~| w794;
assign w877 = w263 ~| w795;
assign w878 = w292 ~| w795;
assign w879 = w243 ~| w796;
assign w880 = w268 ~| w796;
assign w881 = w325 ~| w797;
assign w882 = w233 ~| w797;
assign w883 = w398 ~| w798;
assign w884 = w289 ~| w798;
assign w885 = w313 ~| w800;
assign w886 = w360 ~| w800;
assign w887 = w227 ~| w801;
assign w888 = w348 ~| w801;
assign w889 = ~w808;
assign w890 = w803 ~| w809;
assign w891 = w383 | w818;
assign w892 = w812 ~| w819;
assign w893 = w228 ~| w820;
assign w894 = w309 ~| w820;
assign w895 = w218 ~| w820;
assign w896 = w265 ~| w821;
assign w897 = w389 ~| w821;
assign w898 = w277 ~| w822;
assign w899 = w280 ~| w822;
assign w900 = w325 ~| w823;
assign w901 = w301 ~| w823;
assign w902 = w246 ~| w824;
assign w903 = w338 ~| w824;
assign w904 = w364 ~| w826;
assign w905 = w378 ~| w826;
assign w906 = w257 ~| w827;
assign w907 = w343 ~| w827;
assign w908 = w588 & w829;
assign w909 = w767 | w834;
assign w910 = w304 ~| w837;
assign w911 = w237 ~| w837;
assign w912 = w334 ~| w837;
assign w913 = w265 ~| w838;
assign w914 = w394 ~| w838;
assign w915 = w301 ~| w839;
assign w916 = w321 ~| w839;
assign w917 = w289 ~| w840;
assign w918 = w253 ~| w840;
assign w919 = w245 ~| w841;
assign w920 = w352 ~| w841;
assign w921 = w364 ~| w843;
assign w922 = w277 ~| w843;
assign w923 = w378 ~| w844;
assign w924 = w223 ~| w844;
assign w925 = w152 | w845;
assign w926 = ~w846;
assign w927 = w55 ~^ w848;
assign w928 = w715 | w849;
assign w929 = w485 | w851;
assign w930 = w648 | w853;
assign w931 = w290 ~^ w854;
assign w932 = w291 | w854;
assign w933 = w708 | w855;
assign out1[1] = w708 ^ w855;
assign w934 = w184 ~^ w857;
assign w935 = w709 | w858;
assign w936 = w606 | w859;
assign w937 = w601 | w860;
assign w938 = w598 | w861;
assign w939 = w593 | w863;
assign w940 = w594 | w864;
assign w941 = w597 | w865;
assign w942 = w592 | w866;
assign w943 = w596 | w867;
assign w944 = w600 | w869;
assign w945 = w603 | w870;
assign w946 = w602 | w871;
assign w947 = w599 | w873;
assign w948 = w850 | w874;
assign w949 = w635 | w875;
assign w950 = w739 | w876;
assign w951 = w640 | w878;
assign w952 = w631 | w880;
assign w953 = w630 | w881;
assign w954 = w734 | w883;
assign w955 = w637 | w884;
assign w956 = w634 | w885;
assign w957 = w636 | w886;
assign w958 = w627 | w888;
assign w959 = w657 ~| w889;
assign w960 = w665 & w889;
assign w961 = w187 ~^ w890;
assign w962 = w196 ~^ w891;
assign w963 = w195 ~^ w892;
assign w964 = w746 | w893;
assign w965 = w613 | w894;
assign w966 = w817 | w896;
assign w967 = w619 | w897;
assign w968 = w610 | w899;
assign w969 = w623 | w900;
assign w970 = w852 | w903;
assign w971 = w615 | w904;
assign w972 = w611 | w905;
assign w973 = w614 | w906;
assign w974 = w622 | w907;
assign w975 = w674 | w908;
assign w976 = w586 ~^ w909;
assign w977 = w654 | w910;
assign w978 = w537 | w912;
assign w979 = w644 | w913;
assign w980 = w655 | w917;
assign w981 = w647 | w918;
assign w982 = w656 | w923;
assign w983 = w535 | w924;
assign w984 = w847 ~^ w925;
assign w985 = ~w925;
assign w986 = w846 ~^ w927;
assign w987 = w926 ~| w927;
assign w988 = ~w927;
assign w989 = w554 ~| w929;
assign w990 = w541 ~| w931;
assign w991 = w724 ~| w931;
assign w992 = w497 ~| w931;
assign w993 = w742 ~| w931;
assign w994 = w758 ~| w931;
assign w995 = w437 & w932;
assign w996 = ~w934;
assign w997 = w108 ^ w934;
assign w998 = w114 ~^ w935;
assign w999 = w856 ~| w940;
assign w1000 = w928 ~| w942;
assign w1001 = w804 ~| w948;
assign w1002 = w877 | w959;
assign w1003 = w380 | w960;
assign w1004 = ~w962;
assign w1005 = w136 ^ w962;
assign w1006 = w814 ~| w966;
assign w1007 = w816 ~| w970;
assign w1008 = w584 ~^ w975;
assign w1009 = w682 | w975;
assign w1010 = w682 & w975;
assign w1011 = w930 ~| w978;
assign w1012 = w775 ~| w979;
assign w1013 = ~w984;
assign w1014 = w847 & w985;
assign w1015 = w846 | w988;
assign w1016 = w55 ~^ w989;
assign w1017 = w643 | w990;
assign w1018 = w713 | w991;
assign w1019 = w492 | w992;
assign w1020 = w887 | w993;
assign w1021 = w895 | w994;
assign w1022 = w387 ~^ w995;
assign w1023 = w386 | w995;
assign w1024 = w117 | w996;
assign w1025 = ~w997;
assign w1026 = w113 ^ w999;
assign w1027 = w109 ^ w1000;
assign w1028 = w123 ^ w1001;
assign w1029 = w806 ~| w1002;
assign w1030 = w192 ~^ w1003;
assign w1031 = w141 | w1004;
assign w1032 = ~w1005;
assign w1033 = w197 ~^ w1006;
assign w1034 = w194 ~^ w1007;
assign w1035 = w144 ^ w1011;
assign w1036 = w147 ^ w1012;
assign w1037 = ~w1014;
assign w1038 = w984 ~| w1016;
assign w1039 = ~w1016;
assign w1040 = w983 ~| w1017;
assign w1041 = w936 ~| w1018;
assign w1042 = w551 ~| w1019;
assign w1043 = w802 ~| w1020;
assign w1044 = w815 ~| w1021;
assign w1045 = w541 ~| w1022;
assign w1046 = w758 ~| w1022;
assign w1047 = w497 ~| w1022;
assign w1048 = w724 ~| w1022;
assign w1049 = w742 ~| w1022;
assign w1050 = w463 & w1023;
assign w1051 = ~w1024;
assign w1052 = w998 ^ w1024;
assign w1053 = ~w1026;
assign w1054 = ~w1028;
assign w1055 = w128 ^ w1029;
assign w1056 = ~w1030;
assign w1057 = w127 ^ w1030;
assign w1058 = w963 ~^ w1031;
assign w1059 = ~w1031;
assign w1060 = w574 ~^ w1033;
assign w1061 = w507 ~| w1033;
assign w1062 = ~w1033;
assign w1063 = w576 ~^ w1034;
assign w1064 = w576 ~| w1034;
assign w1065 = w576 & w1034;
assign w1066 = ~w1035;
assign w1067 = w1025 ~| w1036;
assign w1068 = ~w1036;
assign w1069 = w984 ~^ w1039;
assign w1070 = w1013 | w1039;
assign w1071 = w205 ~^ w1040;
assign w1072 = w183 ~^ w1041;
assign w1073 = w106 ^ w1042;
assign w1074 = w126 ^ w1043;
assign w1075 = w198 ~^ w1044;
assign w1076 = w922 | w1045;
assign w1077 = w898 | w1046;
assign w1078 = w491 | w1047;
assign w1079 = w721 | w1048;
assign w1080 = w735 | w1049;
assign w1081 = w388 ~^ w1050;
assign w1082 = w385 | w1050;
assign w1083 = w998 & w1051;
assign w1084 = w1035 ~^ w1052;
assign w1085 = ~w1052;
assign w1086 = w1005 ~^ w1055;
assign w1087 = w1032 ~| w1055;
assign w1088 = ~w1055;
assign w1089 = w129 | w1056;
assign w1090 = w1026 ~^ w1057;
assign w1091 = w1053 | w1057;
assign w1092 = ~w1057;
assign w1093 = w1028 ~^ w1058;
assign w1094 = w1028 ~| w1058;
assign w1095 = ~w1058;
assign w1096 = w963 & w1059;
assign w1097 = w574 | w1062;
assign w1098 = w1052 | w1066;
assign w1099 = w997 | w1068;
assign w1100 = ~w1071;
assign w1101 = ~w1072;
assign w1102 = ~w1073;
assign w1103 = ~w1074;
assign w1104 = w577 ~^ w1075;
assign w1105 = w577 & w1075;
assign w1106 = w577 | w1075;
assign w1107 = w696 ~| w1076;
assign w1108 = w813 ~| w1077;
assign w1109 = w552 ~| w1078;
assign w1110 = w937 ~| w1079;
assign w1111 = w952 ~| w1080;
assign w1112 = w758 ~| w1081;
assign w1113 = w541 ~| w1081;
assign w1114 = w724 ~| w1081;
assign w1115 = w497 ~| w1081;
assign w1116 = w742 ~| w1081;
assign w1117 = w465 & w1082;
assign w1118 = ~w1083;
assign w1119 = w1035 ~| w1085;
assign w1120 = w1005 | w1088;
assign w1121 = w961 ~^ w1089;
assign w1122 = ~w1089;
assign w1123 = w1026 ~| w1092;
assign w1124 = w1054 | w1095;
assign w1125 = ~w1096;
assign w1126 = w145 ^ w1107;
assign w1127 = w63 ~^ w1108;
assign w1128 = w177 ~^ w1109;
assign w1129 = w110 ^ w1110;
assign w1130 = w188 ~^ w1111;
assign w1131 = w901 | w1112;
assign w1132 = w915 | w1113;
assign w1133 = w711 | w1114;
assign w1134 = w484 | w1115;
assign w1135 = w731 | w1116;
assign w1136 = w315 ~^ w1117;
assign w1137 = w314 | w1117;
assign w1138 = w1027 ~^ w1121;
assign w1139 = w1027 & w1121;
assign w1140 = w1027 ~| w1121;
assign w1141 = w961 & w1122;
assign w1142 = ~w1126;
assign w1143 = w688 ~^ w1127;
assign w1144 = w690 & w1127;
assign w1145 = ~w1129;
assign w1146 = ~w1130;
assign w1147 = w811 ~| w1131;
assign w1148 = w698 ~| w1132;
assign w1149 = w946 ~| w1133;
assign w1150 = w547 ~| w1134;
assign w1151 = w951 ~| w1135;
assign w1152 = w758 ~| w1136;
assign w1153 = w541 ~| w1136;
assign w1154 = ~w1136;
assign w1155 = w442 & w1137;
assign w1156 = ~w1141;
assign w1157 = w689 | w1144;
assign w1158 = w196 ~^ w1147;
assign w1159 = w204 ~^ w1148;
assign w1160 = w181 ~^ w1149;
assign w1161 = w55 ~^ w1150;
assign w1162 = w191 ~^ w1151;
assign w1163 = w750 | w1152;
assign w1164 = w914 | w1153;
assign w1165 = ~w1154;
assign w1166 = w808 & w1154;
assign w1167 = w341 ~^ w1155;
assign w1168 = w339 | w1155;
assign w1169 = w683 ~^ w1158;
assign w1170 = w685 & w1158;
assign w1171 = ~w1159;
assign w1172 = ~w1160;
assign w1173 = ~w1162;
assign w1174 = w967 ~| w1163;
assign w1175 = w703 ~| w1164;
assign w1176 = w724 ~| w1165;
assign w1177 = w497 ~| w1165;
assign w1178 = w639 | w1166;
assign w1179 = w742 ~| w1167;
assign w1180 = w497 ~| w1167;
assign w1181 = w724 ~| w1167;
assign w1182 = w541 ~| w1167;
assign w1183 = w758 ~| w1167;
assign w1184 = w451 & w1168;
assign w1185 = w1157 ~^ w1169;
assign w1186 = w1157 & w1169;
assign w1187 = w1157 | w1169;
assign w1188 = w684 | w1170;
assign w1189 = w134 ^ w1174;
assign w1190 = w65 ~^ w1175;
assign w1191 = w719 | w1176;
assign w1192 = w496 | w1177;
assign w1193 = w954 ~| w1178;
assign w1194 = w727 | w1179;
assign w1195 = w494 | w1180;
assign w1196 = w718 | w1181;
assign w1197 = w916 | w1182;
assign w1198 = w757 | w1183;
assign w1199 = w342 ~^ w1184;
assign w1200 = w340 | w1184;
assign w1201 = w670 ~^ w1189;
assign w1202 = w671 & w1189;
assign w1203 = ~w1190;
assign w1204 = w943 ~| w1191;
assign w1205 = w561 ~| w1192;
assign w1206 = w186 ~^ w1193;
assign w1207 = w953 ~| w1194;
assign w1208 = w559 ~| w1195;
assign w1209 = w939 ~| w1196;
assign w1210 = w700 ~| w1197;
assign w1211 = w969 ~| w1198;
assign w1212 = w742 ~| w1199;
assign w1213 = w541 ~| w1199;
assign w1214 = w758 ~| w1199;
assign w1215 = w724 ~| w1199;
assign w1216 = w497 ~| w1199;
assign w1217 = w449 & w1200;
assign w1218 = w1188 ~^ w1201;
assign w1219 = w1188 & w1201;
assign w1220 = w1188 | w1201;
assign w1221 = w672 | w1202;
assign w1222 = w57 ~^ w1204;
assign w1223 = w55 ~^ w1205;
assign w1224 = w61 ~^ w1207;
assign w1225 = w55 ~^ w1208;
assign w1226 = w179 ~^ w1209;
assign w1227 = w202 ~^ w1210;
assign w1228 = w198 ~^ w1211;
assign w1229 = w882 | w1212;
assign w1230 = w911 | w1213;
assign w1231 = w616 | w1214;
assign w1232 = w712 | w1215;
assign w1233 = w489 | w1216;
assign w1234 = w302 ~^ w1217;
assign w1235 = w303 | w1217;
assign w1236 = ~w1223;
assign w1237 = ~w1225;
assign w1238 = ~w1227;
assign w1239 = w675 ~^ w1228;
assign w1240 = w675 & w1228;
assign w1241 = w675 | w1228;
assign w1242 = w805 ~| w1229;
assign w1243 = w697 ~| w1230;
assign w1244 = w964 ~| w1231;
assign w1245 = w944 ~| w1232;
assign w1246 = w558 ~| w1233;
assign w1247 = w742 ~| w1234;
assign w1248 = w497 ~| w1234;
assign w1249 = w724 ~| w1234;
assign w1250 = w541 ~| w1234;
assign w1251 = w758 ~| w1234;
assign w1252 = w439 & w1235;
assign w1253 = w1221 ~^ w1239;
assign w1254 = w1221 & w1241;
assign w1255 = w188 ~^ w1242;
assign w1256 = w65 ~^ w1243;
assign w1257 = w63 ~^ w1244;
assign w1258 = w182 ~^ w1245;
assign w1259 = w55 ~^ w1246;
assign w1260 = w732 | w1247;
assign w1261 = w495 | w1248;
assign w1262 = w710 | w1249;
assign w1263 = w920 | w1250;
assign w1264 = w748 | w1251;
assign w1265 = w278 ~^ w1252;
assign w1266 = w279 | w1252;
assign w1267 = w1240 | w1254;
assign w1268 = w1185 ~^ w1255;
assign w1269 = w1187 & w1255;
assign w1270 = ~w1256;
assign w1271 = w830 ~^ w1257;
assign w1272 = w831 & w1257;
assign w1273 = ~w1259;
assign w1274 = w958 ~| w1260;
assign w1275 = w560 ~| w1261;
assign w1276 = w945 ~| w1262;
assign w1277 = w702 ~| w1263;
assign w1278 = w974 ~| w1264;
assign w1279 = w742 ~| w1265;
assign w1280 = w497 ~| w1265;
assign w1281 = w758 ~| w1265;
assign w1282 = w724 ~| w1265;
assign w1283 = w541 ~| w1265;
assign w1284 = w434 & w1266;
assign w1285 = w1186 | w1269;
assign w1286 = w1267 ~^ w1271;
assign w1287 = ~w1271;
assign w1288 = w832 | w1272;
assign w1289 = w191 ~^ w1274;
assign w1290 = w55 ~^ w1275;
assign w1291 = w184 ~^ w1276;
assign w1292 = w206 ~^ w1277;
assign w1293 = w195 ~^ w1278;
assign w1294 = w738 | w1279;
assign w1295 = w483 | w1280;
assign w1296 = w747 | w1281;
assign w1297 = w872 | w1282;
assign w1298 = w540 | w1283;
assign w1299 = w354 ~^ w1284;
assign w1300 = w353 | w1284;
assign w1301 = w1267 | w1287;
assign w1302 = w1267 & w1287;
assign w1303 = ~w1288;
assign w1304 = w1218 ~^ w1289;
assign w1305 = w1220 & w1289;
assign w1306 = w828 ~^ w1293;
assign w1307 = w760 & w1293;
assign w1308 = w956 ~| w1294;
assign w1309 = w555 ~| w1295;
assign w1310 = w965 ~| w1296;
assign w1311 = w782 ~| w1297;
assign w1312 = w977 ~| w1298;
assign w1313 = w758 ~| w1299;
assign w1314 = w497 ~| w1299;
assign w1315 = w724 ~| w1299;
assign w1316 = w742 ~| w1299;
assign w1317 = w541 ~| w1299;
assign w1318 = w453 & w1300;
assign w1319 = w1285 ~^ w1304;
assign w1320 = w1285 & w1304;
assign w1321 = w1285 | w1304;
assign w1322 = w1219 | w1305;
assign w1323 = w1288 ~^ w1306;
assign w1324 = w1303 ~| w1306;
assign w1325 = ~w1306;
assign w1326 = w763 | w1307;
assign w1327 = w186 ~^ w1308;
assign w1328 = w55 ~^ w1309;
assign w1329 = w199 ~^ w1310;
assign w1330 = w179 ~^ w1311;
assign w1331 = w202 ~^ w1312;
assign w1332 = w749 | w1313;
assign w1333 = w486 | w1314;
assign w1334 = w868 | w1315;
assign w1335 = w629 | w1316;
assign w1336 = w529 | w1317;
assign w1337 = w367 ~^ w1318;
assign w1338 = w365 | w1318;
assign w1339 = w1288 | w1325;
assign w1340 = w1253 ~^ w1327;
assign w1341 = w1253 & w1327;
assign w1342 = w1253 | w1327;
assign w1343 = w770 ~^ w1329;
assign w1344 = w835 | w1329;
assign w1345 = ~w1329;
assign w1346 = w973 ~| w1332;
assign w1347 = w556 ~| w1333;
assign w1348 = w780 ~| w1334;
assign w1349 = w950 ~| w1335;
assign w1350 = w981 ~| w1336;
assign w1351 = w724 ~| w1337;
assign w1352 = w541 ~| w1337;
assign w1353 = w758 ~| w1337;
assign w1354 = w497 ~| w1337;
assign w1355 = w742 ~| w1337;
assign w1356 = w458 & w1338;
assign w1357 = w1322 ~^ w1340;
assign w1358 = w1322 & w1342;
assign w1359 = w1326 ~^ w1343;
assign w1360 = w1326 & w1344;
assign w1361 = w770 ~| w1345;
assign w1362 = w63 ~^ w1346;
assign w1363 = w55 ~^ w1347;
assign w1364 = w112 ^ w1348;
assign w1365 = w61 ~^ w1349;
assign w1366 = w146 ^ w1350;
assign w1367 = w716 | w1351;
assign w1368 = w539 | w1352;
assign w1369 = w753 | w1353;
assign w1370 = w487 | w1354;
assign w1371 = w733 | w1355;
assign w1372 = w368 ~^ w1356;
assign w1373 = w366 | w1356;
assign w1374 = w1341 | w1358;
assign w1375 = ~w1359;
assign w1376 = w1360 | w1361;
assign w1377 = w1008 ~^ w1362;
assign w1378 = w1009 & w1362;
assign w1379 = w1286 ~^ w1365;
assign w1380 = w1301 & w1365;
assign w1381 = w938 ~| w1367;
assign w1382 = w980 ~| w1368;
assign w1383 = w968 ~| w1369;
assign w1384 = w549 ~| w1370;
assign w1385 = w955 ~| w1371;
assign w1386 = w497 ~| w1372;
assign w1387 = w742 ~| w1372;
assign w1388 = w724 ~| w1372;
assign w1389 = w541 ~| w1372;
assign w1390 = w758 ~| w1372;
assign w1391 = w456 & w1373;
assign w1392 = ~w1374;
assign w1393 = ~w1376;
assign w1394 = w1376 ~^ w1377;
assign w1395 = ~w1377;
assign w1396 = w1010 | w1378;
assign w1397 = w1374 ~^ w1379;
assign w1398 = ~w1379;
assign w1399 = w1302 | w1380;
assign w1400 = w57 ~^ w1381;
assign w1401 = w65 ~^ w1382;
assign w1402 = w199 ~^ w1383;
assign w1403 = w55 ~^ w1384;
assign w1404 = w190 ~^ w1385;
assign w1405 = w490 | w1386;
assign w1406 = w729 | w1387;
assign w1407 = w717 | w1388;
assign w1408 = w921 | w1389;
assign w1409 = w755 | w1390;
assign w1410 = w247 | w1391;
assign w1411 = ~w1391;
assign w1412 = w1379 ~| w1392;
assign w1413 = w1377 ~| w1393;
assign w1414 = w1376 | w1395;
assign w1415 = ~w1396;
assign w1416 = w1374 | w1398;
assign w1417 = ~w1399;
assign w1418 = w1319 ~^ w1400;
assign w1419 = w1321 & w1400;
assign w1420 = w833 ~^ w1402;
assign w1421 = w765 & w1402;
assign w1422 = w1323 ~^ w1404;
assign w1423 = w1339 & w1404;
assign w1424 = w550 ~| w1405;
assign w1425 = w957 ~| w1406;
assign w1426 = w941 ~| w1407;
assign w1427 = w701 ~| w1408;
assign w1428 = w971 ~| w1409;
assign w1429 = w758 ~| w1410;
assign w1430 = ~w1410;
assign w1431 = w497 ~| w1410;
assign w1432 = w724 ~| w1410;
assign w1433 = w541 ~| w1410;
assign w1434 = w161 ~| w1411;
assign w1435 = ~w1418;
assign w1436 = w1320 | w1419;
assign w1437 = w1396 ~^ w1420;
assign w1438 = w768 | w1421;
assign w1439 = w1399 ~^ w1422;
assign w1440 = w1324 | w1423;
assign w1441 = w55 ~^ w1424;
assign w1442 = w189 ~^ w1425;
assign w1443 = w180 ~^ w1426;
assign w1444 = w203 ~^ w1427;
assign w1445 = w63 ~^ w1428;
assign w1446 = w902 | w1429;
assign w1447 = ~w1430;
assign w1448 = w481 | w1431;
assign w1449 = w862 | w1432;
assign w1450 = w919 | w1433;
assign w1451 = w1430 | w1434;
assign w1452 = w1359 ~^ w1442;
assign w1453 = w1375 | w1442;
assign w1454 = ~w1442;
assign w1455 = w1357 ~^ w1443;
assign w1456 = w1357 & w1443;
assign w1457 = w1357 | w1443;
assign w1458 = ~w1444;
assign w1459 = w771 ~^ w1445;
assign w1460 = w836 | w1445;
assign w1461 = ~w1445;
assign w1462 = w137 ^ w1446;
assign w1463 = w742 ~| w1447;
assign w1464 = w55 ~^ w1448;
assign w1465 = w57 ~^ w1449;
assign w1466 = w65 ~^ w1450;
assign w1467 = w541 ~| w1451;
assign w1468 = w758 ~| w1451;
assign w1469 = w497 ~| w1451;
assign w1470 = w724 ~| w1451;
assign w1471 = w742 ~| w1451;
assign w1472 = w1440 ~^ w1452;
assign w1473 = w1440 & w1453;
assign w1474 = w1359 ~| w1454;
assign w1475 = w1436 ~^ w1455;
assign w1476 = w1436 & w1457;
assign w1477 = w1438 ~^ w1459;
assign w1478 = w1438 & w1460;
assign w1479 = w771 ~| w1461;
assign w1480 = w686 ~^ w1462;
assign w1481 = w879 | w1463;
assign w1482 = ~w1464;
assign w1483 = w1439 ~^ w1465;
assign w1484 = w1417 | w1465;
assign w1485 = ~w1465;
assign w1486 = w982 ~| w1467;
assign w1487 = w972 ~| w1468;
assign w1488 = w553 ~| w1469;
assign w1489 = w947 ~| w1470;
assign w1490 = w949 ~| w1471;
assign w1491 = w1473 | w1474;
assign w1492 = ~w1475;
assign w1493 = w1456 | w1476;
assign w1494 = w1478 | w1479;
assign w1495 = w124 ^ w1481;
assign w1496 = w1399 ~| w1485;
assign w1497 = w205 ~^ w1486;
assign w1498 = w138 ^ w1487;
assign w1499 = w55 ~^ w1488;
assign w1500 = w57 ~^ w1489;
assign w1501 = w189 ~^ w1490;
assign w1502 = ~w1491;
assign w1503 = ~w1493;
assign w1504 = ~w1494;
assign w1505 = w1437 ~^ w1495;
assign w1506 = w1415 | w1495;
assign w1507 = ~w1495;
assign w1508 = w1422 | w1496;
assign w1509 = w976 ~^ w1498;
assign w1510 = w1397 ~^ w1500;
assign w1511 = w1416 & w1500;
assign w1512 = w1394 ~^ w1501;
assign w1513 = w1414 & w1501;
assign w1514 = w1396 ~| w1507;
assign w1515 = w1484 & w1508;
assign w1516 = w1494 ~^ w1509;
assign w1517 = w1504 ~| w1509;
assign w1518 = w1504 & w1509;
assign w1519 = w1493 ~^ w1510;
assign w1520 = w1503 ~| w1510;
assign w1521 = w1503 & w1510;
assign w1522 = w1412 | w1511;
assign w1523 = w1491 ~^ w1512;
assign w1524 = w1502 ~| w1512;
assign w1525 = w1502 & w1512;
assign w1526 = w1413 | w1513;
assign w1527 = w1420 | w1514;
assign w1528 = w1472 ~^ w1515;
assign w1529 = w1472 & w1515;
assign w1530 = w1472 | w1515;
assign w1531 = w1483 ~^ w1522;
assign w1532 = w1483 & w1522;
assign w1533 = w1483 | w1522;
assign w1534 = w1505 ~^ w1526;
assign w1535 = w1505 & w1526;
assign w1536 = w1505 | w1526;
assign w1537 = w1506 & w1527;
assign w1538 = w1477 ~^ w1537;
assign w1539 = w1477 | w1537;
assign w1540 = w1477 & w1537;
wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540;
endmodule